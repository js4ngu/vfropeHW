module Int64ToFP32(
  input  [63:0] io_inInt,
  output [31:0] io_outIEEE
);
  wire  sign = io_inInt[63]; // @[FPU.scala 139:22]
  wire [63:0] _absVal_T_5 = 64'sh0 - $signed(io_inInt); // @[FPU.scala 140:79]
  wire [63:0] _absVal_T_7 = sign ? _absVal_T_5 : io_inInt; // @[FPU.scala 140:46]
  wire [63:0] absVal = $signed(io_inInt) == 64'sh0 ? 64'h0 : _absVal_T_7; // @[FPU.scala 140:19]
  wire  isZero = absVal == 64'h0; // @[FPU.scala 141:23]
  wire [63:0] _GEN_0 = {{32'd0}, absVal[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_3 = _GEN_0 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_5 = {absVal[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_7 = _LeadingOne_T_5 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_8 = _LeadingOne_T_3 | _LeadingOne_T_7; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_1 = {{16'd0}, _LeadingOne_T_8[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_13 = _GEN_1 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_15 = {_LeadingOne_T_8[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_17 = _LeadingOne_T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_18 = _LeadingOne_T_13 | _LeadingOne_T_17; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_2 = {{8'd0}, _LeadingOne_T_18[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_23 = _GEN_2 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_25 = {_LeadingOne_T_18[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_27 = _LeadingOne_T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_28 = _LeadingOne_T_23 | _LeadingOne_T_27; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_3 = {{4'd0}, _LeadingOne_T_28[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_33 = _GEN_3 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_35 = {_LeadingOne_T_28[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_37 = _LeadingOne_T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_38 = _LeadingOne_T_33 | _LeadingOne_T_37; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_4 = {{2'd0}, _LeadingOne_T_38[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_43 = _GEN_4 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_45 = {_LeadingOne_T_38[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_47 = _LeadingOne_T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_48 = _LeadingOne_T_43 | _LeadingOne_T_47; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_5 = {{1'd0}, _LeadingOne_T_48[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_53 = _GEN_5 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _LeadingOne_T_55 = {_LeadingOne_T_48[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _LeadingOne_T_57 = _LeadingOne_T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] _LeadingOne_T_58 = _LeadingOne_T_53 | _LeadingOne_T_57; // @[Bitwise.scala 108:39]
  wire [5:0] _LeadingOne_T_123 = _LeadingOne_T_58[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_124 = _LeadingOne_T_58[61] ? 6'h3d : _LeadingOne_T_123; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_125 = _LeadingOne_T_58[60] ? 6'h3c : _LeadingOne_T_124; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_126 = _LeadingOne_T_58[59] ? 6'h3b : _LeadingOne_T_125; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_127 = _LeadingOne_T_58[58] ? 6'h3a : _LeadingOne_T_126; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_128 = _LeadingOne_T_58[57] ? 6'h39 : _LeadingOne_T_127; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_129 = _LeadingOne_T_58[56] ? 6'h38 : _LeadingOne_T_128; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_130 = _LeadingOne_T_58[55] ? 6'h37 : _LeadingOne_T_129; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_131 = _LeadingOne_T_58[54] ? 6'h36 : _LeadingOne_T_130; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_132 = _LeadingOne_T_58[53] ? 6'h35 : _LeadingOne_T_131; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_133 = _LeadingOne_T_58[52] ? 6'h34 : _LeadingOne_T_132; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_134 = _LeadingOne_T_58[51] ? 6'h33 : _LeadingOne_T_133; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_135 = _LeadingOne_T_58[50] ? 6'h32 : _LeadingOne_T_134; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_136 = _LeadingOne_T_58[49] ? 6'h31 : _LeadingOne_T_135; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_137 = _LeadingOne_T_58[48] ? 6'h30 : _LeadingOne_T_136; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_138 = _LeadingOne_T_58[47] ? 6'h2f : _LeadingOne_T_137; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_139 = _LeadingOne_T_58[46] ? 6'h2e : _LeadingOne_T_138; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_140 = _LeadingOne_T_58[45] ? 6'h2d : _LeadingOne_T_139; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_141 = _LeadingOne_T_58[44] ? 6'h2c : _LeadingOne_T_140; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_142 = _LeadingOne_T_58[43] ? 6'h2b : _LeadingOne_T_141; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_143 = _LeadingOne_T_58[42] ? 6'h2a : _LeadingOne_T_142; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_144 = _LeadingOne_T_58[41] ? 6'h29 : _LeadingOne_T_143; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_145 = _LeadingOne_T_58[40] ? 6'h28 : _LeadingOne_T_144; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_146 = _LeadingOne_T_58[39] ? 6'h27 : _LeadingOne_T_145; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_147 = _LeadingOne_T_58[38] ? 6'h26 : _LeadingOne_T_146; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_148 = _LeadingOne_T_58[37] ? 6'h25 : _LeadingOne_T_147; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_149 = _LeadingOne_T_58[36] ? 6'h24 : _LeadingOne_T_148; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_150 = _LeadingOne_T_58[35] ? 6'h23 : _LeadingOne_T_149; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_151 = _LeadingOne_T_58[34] ? 6'h22 : _LeadingOne_T_150; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_152 = _LeadingOne_T_58[33] ? 6'h21 : _LeadingOne_T_151; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_153 = _LeadingOne_T_58[32] ? 6'h20 : _LeadingOne_T_152; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_154 = _LeadingOne_T_58[31] ? 6'h1f : _LeadingOne_T_153; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_155 = _LeadingOne_T_58[30] ? 6'h1e : _LeadingOne_T_154; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_156 = _LeadingOne_T_58[29] ? 6'h1d : _LeadingOne_T_155; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_157 = _LeadingOne_T_58[28] ? 6'h1c : _LeadingOne_T_156; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_158 = _LeadingOne_T_58[27] ? 6'h1b : _LeadingOne_T_157; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_159 = _LeadingOne_T_58[26] ? 6'h1a : _LeadingOne_T_158; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_160 = _LeadingOne_T_58[25] ? 6'h19 : _LeadingOne_T_159; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_161 = _LeadingOne_T_58[24] ? 6'h18 : _LeadingOne_T_160; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_162 = _LeadingOne_T_58[23] ? 6'h17 : _LeadingOne_T_161; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_163 = _LeadingOne_T_58[22] ? 6'h16 : _LeadingOne_T_162; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_164 = _LeadingOne_T_58[21] ? 6'h15 : _LeadingOne_T_163; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_165 = _LeadingOne_T_58[20] ? 6'h14 : _LeadingOne_T_164; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_166 = _LeadingOne_T_58[19] ? 6'h13 : _LeadingOne_T_165; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_167 = _LeadingOne_T_58[18] ? 6'h12 : _LeadingOne_T_166; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_168 = _LeadingOne_T_58[17] ? 6'h11 : _LeadingOne_T_167; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_169 = _LeadingOne_T_58[16] ? 6'h10 : _LeadingOne_T_168; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_170 = _LeadingOne_T_58[15] ? 6'hf : _LeadingOne_T_169; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_171 = _LeadingOne_T_58[14] ? 6'he : _LeadingOne_T_170; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_172 = _LeadingOne_T_58[13] ? 6'hd : _LeadingOne_T_171; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_173 = _LeadingOne_T_58[12] ? 6'hc : _LeadingOne_T_172; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_174 = _LeadingOne_T_58[11] ? 6'hb : _LeadingOne_T_173; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_175 = _LeadingOne_T_58[10] ? 6'ha : _LeadingOne_T_174; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_176 = _LeadingOne_T_58[9] ? 6'h9 : _LeadingOne_T_175; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_177 = _LeadingOne_T_58[8] ? 6'h8 : _LeadingOne_T_176; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_178 = _LeadingOne_T_58[7] ? 6'h7 : _LeadingOne_T_177; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_179 = _LeadingOne_T_58[6] ? 6'h6 : _LeadingOne_T_178; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_180 = _LeadingOne_T_58[5] ? 6'h5 : _LeadingOne_T_179; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_181 = _LeadingOne_T_58[4] ? 6'h4 : _LeadingOne_T_180; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_182 = _LeadingOne_T_58[3] ? 6'h3 : _LeadingOne_T_181; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_183 = _LeadingOne_T_58[2] ? 6'h2 : _LeadingOne_T_182; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_184 = _LeadingOne_T_58[1] ? 6'h1 : _LeadingOne_T_183; // @[Mux.scala 47:70]
  wire [5:0] _LeadingOne_T_185 = _LeadingOne_T_58[0] ? 6'h0 : _LeadingOne_T_184; // @[Mux.scala 47:70]
  wire [5:0] LeadingOne = isZero ? 6'h0 : _LeadingOne_T_185; // @[FPU.scala 144:23]
  wire [5:0] shiftAmount = isZero ? 6'h0 : LeadingOne; // @[FPU.scala 147:24]
  wire [126:0] _GEN_7 = {{63'd0}, absVal}; // @[FPU.scala 148:53]
  wire [126:0] _normalizedMantissa_T = _GEN_7 << shiftAmount; // @[FPU.scala 148:53]
  wire [22:0] normalizedMantissa = isZero ? 23'h0 : _normalizedMantissa_T[62:40]; // @[FPU.scala 148:31]
  wire [7:0] _GEN_6 = {{2'd0}, LeadingOne}; // @[FPU.scala 151:48]
  wire [7:0] _biasedExponent_T_1 = 8'hbe - _GEN_6; // @[FPU.scala 151:48]
  wire [7:0] biasedExponent = isZero ? 8'h0 : _biasedExponent_T_1; // @[FPU.scala 151:27]
  wire [8:0] outIEEE_hi = {sign,biasedExponent}; // @[Cat.scala 33:92]
  assign io_outIEEE = {outIEEE_hi,normalizedMantissa}; // @[Cat.scala 33:92]
endmodule
module MulFullRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [47:0] io_rawOut_sig
);
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isZero | io_a_isZero & io_b_isInf; // @[MulRecFN.scala 58:60]
  wire [9:0] _common_sExpOut_T_2 = $signed(io_a_sExp) + $signed(io_b_sExp); // @[MulRecFN.scala 62:36]
  wire [49:0] _common_sigOut_T = io_a_sig * io_b_sig; // @[MulRecFN.scala 63:35]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[MulRecFN.scala 66:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[MulRecFN.scala 70:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[MulRecFN.scala 59:38]
  assign io_rawOut_isZero = io_a_isZero | io_b_isZero; // @[MulRecFN.scala 60:40]
  assign io_rawOut_sign = io_a_sign ^ io_b_sign; // @[MulRecFN.scala 61:36]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - 10'sh100; // @[MulRecFN.scala 62:48]
  assign io_rawOut_sig = _common_sigOut_T[47:0]; // @[MulRecFN.scala 63:46]
endmodule
module MulRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  mulFullRaw_io_a_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_a_sExp; // @[MulRecFN.scala 84:28]
  wire [24:0] mulFullRaw_io_a_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_b_sExp; // @[MulRecFN.scala 84:28]
  wire [24:0] mulFullRaw_io_b_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_invalidExc; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 84:28]
  wire [47:0] mulFullRaw_io_rawOut_sig; // @[MulRecFN.scala 84:28]
  wire  _io_rawOut_sig_T_2 = |mulFullRaw_io_rawOut_sig[21:0]; // @[MulRecFN.scala 93:55]
  MulFullRawFN mulFullRaw ( // @[MulRecFN.scala 84:28]
    .io_a_isNaN(mulFullRaw_io_a_isNaN),
    .io_a_isInf(mulFullRaw_io_a_isInf),
    .io_a_isZero(mulFullRaw_io_a_isZero),
    .io_a_sign(mulFullRaw_io_a_sign),
    .io_a_sExp(mulFullRaw_io_a_sExp),
    .io_a_sig(mulFullRaw_io_a_sig),
    .io_b_isNaN(mulFullRaw_io_b_isNaN),
    .io_b_isInf(mulFullRaw_io_b_isInf),
    .io_b_isZero(mulFullRaw_io_b_isZero),
    .io_b_sign(mulFullRaw_io_b_sign),
    .io_b_sExp(mulFullRaw_io_b_sExp),
    .io_b_sig(mulFullRaw_io_b_sig),
    .io_invalidExc(mulFullRaw_io_invalidExc),
    .io_rawOut_isNaN(mulFullRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(mulFullRaw_io_rawOut_isInf),
    .io_rawOut_isZero(mulFullRaw_io_rawOut_isZero),
    .io_rawOut_sign(mulFullRaw_io_rawOut_sign),
    .io_rawOut_sExp(mulFullRaw_io_rawOut_sExp),
    .io_rawOut_sig(mulFullRaw_io_rawOut_sig)
  );
  assign io_invalidExc = mulFullRaw_io_invalidExc; // @[MulRecFN.scala 89:19]
  assign io_rawOut_isNaN = mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isInf = mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isZero = mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sign = mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sExp = mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sig = {mulFullRaw_io_rawOut_sig[47:22],_io_rawOut_sig_T_2}; // @[Cat.scala 33:92]
  assign mulFullRaw_io_a_isNaN = io_a_isNaN; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isInf = io_a_isInf; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isZero = io_a_isZero; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sign = io_a_sign; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sExp = io_a_sExp; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sig = io_a_sig; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_b_isNaN = io_b_isNaN; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isInf = io_b_isInf; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isZero = io_b_isZero; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sign = io_b_sign; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sExp = io_b_sExp; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sig = io_b_sig; // @[MulRecFN.scala 87:21]
endmodule
module RoundAnyRawFNToRecFN_ie8_is26_oe8_os24(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 120:57]
  wire [8:0] _roundMask_T_1 = ~io_in_sExp[8:0]; // @[primitives.scala 52:21]
  wire  roundMask_msb = _roundMask_T_1[8]; // @[primitives.scala 58:25]
  wire [7:0] roundMask_lsbs = _roundMask_T_1[7:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_1 = roundMask_lsbs[7]; // @[primitives.scala 58:25]
  wire [6:0] roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[6]; // @[primitives.scala 58:25]
  wire [5:0] roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[primitives.scala 59:26]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> roundMask_lsbs_2; // @[primitives.scala 76:56]
  wire [15:0] _GEN_0 = {{8'd0}, roundMask_shift[57:50]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_7 = _GEN_0 & 16'hff; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_9 = {roundMask_shift[49:42], 8'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_11 = _roundMask_T_9 & 16'hff00; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_1 = {{4'd0}, _roundMask_T_12[15:4]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_17 = _GEN_1 & 16'hf0f; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_19 = {_roundMask_T_12[11:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_21 = _roundMask_T_19 & 16'hf0f0; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_2 = {{2'd0}, _roundMask_T_22[15:2]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_27 = _GEN_2 & 16'h3333; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_29 = {_roundMask_T_22[13:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_31 = _roundMask_T_29 & 16'hcccc; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_3 = {{1'd0}, _roundMask_T_32[15:1]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_37 = _GEN_3 & 16'h5555; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_39 = {_roundMask_T_32[14:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_41 = _roundMask_T_39 & 16'haaaa; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 108:39]
  wire [21:0] _roundMask_T_59 = {_roundMask_T_42,roundMask_shift[58],roundMask_shift[59],roundMask_shift[60],
    roundMask_shift[61],roundMask_shift[62],roundMask_shift[63]}; // @[Cat.scala 33:92]
  wire [21:0] _roundMask_T_60 = ~_roundMask_T_59; // @[primitives.scala 73:32]
  wire [21:0] _roundMask_T_61 = roundMask_msb_2 ? 22'h0 : _roundMask_T_60; // @[primitives.scala 73:21]
  wire [21:0] _roundMask_T_62 = ~_roundMask_T_61; // @[primitives.scala 73:17]
  wire [24:0] _roundMask_T_63 = {_roundMask_T_62,3'h7}; // @[primitives.scala 68:58]
  wire [2:0] _roundMask_T_70 = {roundMask_shift[0],roundMask_shift[1],roundMask_shift[2]}; // @[Cat.scala 33:92]
  wire [2:0] _roundMask_T_71 = roundMask_msb_2 ? _roundMask_T_70 : 3'h0; // @[primitives.scala 62:24]
  wire [24:0] _roundMask_T_72 = roundMask_msb_1 ? _roundMask_T_63 : {{22'd0}, _roundMask_T_71}; // @[primitives.scala 67:24]
  wire [24:0] _roundMask_T_73 = roundMask_msb ? _roundMask_T_72 : 25'h0; // @[primitives.scala 62:24]
  wire [24:0] _GEN_4 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [24:0] _roundMask_T_74 = _roundMask_T_73 | _GEN_4; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [26:0] roundMask = {_roundMask_T_74,2'h3}; // @[RoundAnyRawFNToRecFN.scala 159:42]
  wire [27:0] _shiftedRoundMask_T = {1'h0,_roundMask_T_74,2'h3}; // @[RoundAnyRawFNToRecFN.scala 162:41]
  wire [26:0] shiftedRoundMask = _shiftedRoundMask_T[27:1]; // @[RoundAnyRawFNToRecFN.scala 162:53]
  wire [26:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:28]
  wire [26:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 163:46]
  wire [26:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 164:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 164:56]
  wire [26:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 165:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 165:62]
  wire [26:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 174:32]
  wire [25:0] _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 174:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 176:30]
  wire [25:0] _roundedSig_T_7 = roundPosBit & _roundedSig_T_4 ? roundMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 175:25]
  wire [25:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 175:21]
  wire [25:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 174:57]
  wire [26:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 180:32]
  wire [26:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 180:30]
  wire [25:0] _roundedSig_T_16 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 180:47]
  wire [25:0] roundedSig = roundPosBit ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 173:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 185:76]
  wire [9:0] _GEN_5 = {{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [10:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [8:0] common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 187:37]
  wire [22:0] common_fractOut = doShiftSigDown1 ? roundedSig[23:1] : roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:16]
  wire [3:0] _common_overflow_T = sRoundedExp[10:7]; // @[RoundAnyRawFNToRecFN.scala 196:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 196:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 200:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 235:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 237:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 238:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 248:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 250:22]
  wire [8:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 253:18]
  wire [8:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 253:14]
  wire [8:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 252:24]
  wire [8:0] _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 265:18]
  wire [8:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 265:14]
  wire [8:0] _expOut_T_13 = _expOut_T_3 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 264:17]
  wire [8:0] _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 277:16]
  wire [8:0] _expOut_T_19 = _expOut_T_13 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 276:15]
  wire [8:0] _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 278:16]
  wire [8:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 277:73]
  wire [22:0] _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 281:16]
  wire [22:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 280:12]
  wire [9:0] _io_out_T = {signOut,expOut}; // @[RoundAnyRawFNToRecFN.scala 286:23]
  assign io_out = {_io_out_T,fractOut}; // @[RoundAnyRawFNToRecFN.scala 286:33]
endmodule
module RoundRawFNToRecFN_e8_s24(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 310:15]
  RoundAnyRawFNToRecFN_ie8_is26_oe8_os24 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 310:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 318:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 315:44]
endmodule
module MulRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  output [32:0] io_out
);
  wire  mulRawFN__io_a_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_a_sExp; // @[MulRecFN.scala 113:26]
  wire [24:0] mulRawFN__io_a_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_b_sExp; // @[MulRecFN.scala 113:26]
  wire [24:0] mulRawFN__io_b_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_invalidExc; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 113:26]
  wire [26:0] mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 113:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulRecFN.scala 121:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[MulRecFN.scala 121:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[MulRecFN.scala 121:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[MulRecFN.scala 121:15]
  wire [8:0] mulRawFN_io_a_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  mulRawFN_io_a_isZero = mulRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  mulRawFN_io_a_isSpecial = mulRawFN_io_a_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _mulRawFN_io_a_out_sig_T = ~mulRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _mulRawFN_io_a_out_sig_T_1 = {1'h0,_mulRawFN_io_a_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  wire [8:0] mulRawFN_io_b_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  mulRawFN_io_b_isZero = mulRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  mulRawFN_io_b_isSpecial = mulRawFN_io_b_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _mulRawFN_io_b_out_sig_T = ~mulRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _mulRawFN_io_b_out_sig_T_1 = {1'h0,_mulRawFN_io_b_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  MulRawFN mulRawFN_ ( // @[MulRecFN.scala 113:26]
    .io_a_isNaN(mulRawFN__io_a_isNaN),
    .io_a_isInf(mulRawFN__io_a_isInf),
    .io_a_isZero(mulRawFN__io_a_isZero),
    .io_a_sign(mulRawFN__io_a_sign),
    .io_a_sExp(mulRawFN__io_a_sExp),
    .io_a_sig(mulRawFN__io_a_sig),
    .io_b_isNaN(mulRawFN__io_b_isNaN),
    .io_b_isInf(mulRawFN__io_b_isInf),
    .io_b_isZero(mulRawFN__io_b_isZero),
    .io_b_sign(mulRawFN__io_b_sign),
    .io_b_sExp(mulRawFN__io_b_sExp),
    .io_b_sig(mulRawFN__io_b_sig),
    .io_invalidExc(mulRawFN__io_invalidExc),
    .io_rawOut_isNaN(mulRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(mulRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(mulRawFN__io_rawOut_isZero),
    .io_rawOut_sign(mulRawFN__io_rawOut_sign),
    .io_rawOut_sExp(mulRawFN__io_rawOut_sExp),
    .io_rawOut_sig(mulRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN_e8_s24 roundRawFNToRecFN ( // @[MulRecFN.scala 121:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[MulRecFN.scala 127:23]
  assign mulRawFN__io_a_isNaN = mulRawFN_io_a_isSpecial & mulRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_a_isInf = mulRawFN_io_a_isSpecial & ~mulRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign mulRawFN__io_a_isZero = mulRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign mulRawFN__io_a_sign = io_a[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign mulRawFN__io_a_sExp = {1'b0,$signed(mulRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign mulRawFN__io_a_sig = {_mulRawFN_io_a_out_sig_T_1,io_a[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign mulRawFN__io_b_isNaN = mulRawFN_io_b_isSpecial & mulRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_b_isInf = mulRawFN_io_b_isSpecial & ~mulRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign mulRawFN__io_b_isZero = mulRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign mulRawFN__io_b_sign = io_b[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign mulRawFN__io_b_sExp = {1'b0,$signed(mulRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign mulRawFN__io_b_sig = {_mulRawFN_io_b_out_sig_T_1,io_b[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign roundRawFNToRecFN_io_invalidExc = mulRawFN__io_invalidExc; // @[MulRecFN.scala 122:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isInf = mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isZero = mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sign = mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sExp = mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sig = mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 124:39]
endmodule
module FP32Multiplier(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire [32:0] mulRecFN_io_a; // @[FPU.scala 88:26]
  wire [32:0] mulRecFN_io_b; // @[FPU.scala 88:26]
  wire [32:0] mulRecFN_io_out; // @[FPU.scala 88:26]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = mulRecFN_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = mulRecFN_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,mulRecFN_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  MulRecFN mulRecFN ( // @[FPU.scala 88:26]
    .io_a(mulRecFN_io_a),
    .io_b(mulRecFN_io_b),
    .io_out(mulRecFN_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign mulRecFN_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign mulRecFN_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module FP32DivPOW2(
  input  [31:0] io_a,
  output [31:0] io_result
);
  wire [7:0] exponent = io_a[30:23]; // @[FPU.scala 169:22]
  wire [22:0] mantissa = io_a[22:0]; // @[FPU.scala 170:22]
  wire [11:0] _GEN_0 = {{4'd0}, exponent}; // @[FPU.scala 173:30]
  wire [12:0] newExponent = _GEN_0 - 12'h1; // @[FPU.scala 173:30]
  wire  isLessThanZero = newExponent < 13'h7f; // @[FPU.scala 176:36]
  wire [12:0] saturatedExponent = isLessThanZero ? 13'h0 : newExponent; // @[FPU.scala 179:30]
  wire [22:0] saturatedMantissa = isLessThanZero ? 23'h0 : mantissa; // @[FPU.scala 180:30]
  wire [36:0] _io_result_T = {1'h0,saturatedExponent,saturatedMantissa}; // @[Cat.scala 33:92]
  assign io_result = _io_result_T[31:0]; // @[FPU.scala 183:13]
endmodule
module FP32Truncate(
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire  sign = io_in[31]; // @[FPU.scala 195:19]
  wire [7:0] exponent = io_in[30:23]; // @[FPU.scala 196:23]
  wire [22:0] mantissa = io_in[22:0]; // @[FPU.scala 197:23]
  wire [7:0] shift = exponent - 8'h7f; // @[FPU.scala 208:26]
  wire [277:0] _mask_T = 278'h1 << shift; // @[FPU.scala 210:25]
  wire [277:0] _mask_T_2 = _mask_T - 278'h1; // @[FPU.scala 210:35]
  wire [7:0] _mask_T_4 = 8'h17 - shift; // @[FPU.scala 210:51]
  wire [532:0] _GEN_1 = {{255'd0}, _mask_T_2}; // @[FPU.scala 210:42]
  wire [532:0] _mask_T_5 = _GEN_1 << _mask_T_4; // @[FPU.scala 210:42]
  wire [22:0] mask = _mask_T_5[22:0]; // @[FPU.scala 209:20 210:10]
  wire [22:0] truncated_mantissa = mantissa & mask; // @[FPU.scala 212:36]
  wire [31:0] _result_T = {sign,exponent,truncated_mantissa}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_0 = exponent >= 8'h96 ? io_in : _result_T; // @[FPU.scala 203:33 205:12 213:12]
  assign io_out = exponent < 8'h7f ? 32'h0 : _GEN_0; // @[FPU.scala 200:26 202:12]
endmodule
module FP32DivPOW2INT(
  input  [31:0] io_a,
  output [31:0] io_result
);
  wire [31:0] FP32Div_io_a; // @[FPU.scala 225:23]
  wire [31:0] FP32Div_io_result; // @[FPU.scala 225:23]
  wire [31:0] FP32Truncate_io_in; // @[FPU.scala 229:28]
  wire [31:0] FP32Truncate_io_out; // @[FPU.scala 229:28]
  FP32DivPOW2 FP32Div ( // @[FPU.scala 225:23]
    .io_a(FP32Div_io_a),
    .io_result(FP32Div_io_result)
  );
  FP32Truncate FP32Truncate ( // @[FPU.scala 229:28]
    .io_in(FP32Truncate_io_in),
    .io_out(FP32Truncate_io_out)
  );
  assign io_result = FP32Truncate_io_out; // @[FPU.scala 232:13]
  assign FP32Div_io_a = io_a; // @[FPU.scala 226:16]
  assign FP32Truncate_io_in = FP32Div_io_result; // @[FPU.scala 230:22]
endmodule
module AddRawFN(
  input         io_subOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  effSignB = io_b_sign ^ io_subOp; // @[AddRecFN.scala 60:30]
  wire  eqSigns = io_a_sign == effSignB; // @[AddRecFN.scala 61:29]
  wire [9:0] sDiffExps = $signed(io_a_sExp) - $signed(io_b_sExp); // @[AddRecFN.scala 63:31]
  wire  _modNatAlignDist_T = $signed(sDiffExps) < 10'sh0; // @[AddRecFN.scala 64:41]
  wire [9:0] _modNatAlignDist_T_3 = $signed(io_b_sExp) - $signed(io_a_sExp); // @[AddRecFN.scala 64:58]
  wire [9:0] _modNatAlignDist_T_4 = $signed(sDiffExps) < 10'sh0 ? $signed(_modNatAlignDist_T_3) : $signed(sDiffExps); // @[AddRecFN.scala 64:30]
  wire [4:0] modNatAlignDist = _modNatAlignDist_T_4[4:0]; // @[AddRecFN.scala 64:81]
  wire [4:0] _isMaxAlign_T = sDiffExps[9:5]; // @[AddRecFN.scala 66:19]
  wire  _isMaxAlign_T_6 = $signed(_isMaxAlign_T) != -5'sh1 | sDiffExps[4:0] == 5'h0; // @[AddRecFN.scala 67:51]
  wire  isMaxAlign = $signed(_isMaxAlign_T) != 5'sh0 & _isMaxAlign_T_6; // @[AddRecFN.scala 66:45]
  wire [4:0] alignDist = isMaxAlign ? 5'h1f : modNatAlignDist; // @[AddRecFN.scala 68:24]
  wire  _closeSubMags_T = ~eqSigns; // @[AddRecFN.scala 69:24]
  wire  closeSubMags = ~eqSigns & ~isMaxAlign & modNatAlignDist <= 5'h1; // @[AddRecFN.scala 69:48]
  wire  _close_alignedSigA_T = 10'sh0 <= $signed(sDiffExps); // @[AddRecFN.scala 73:18]
  wire [26:0] _close_alignedSigA_T_3 = {io_a_sig, 2'h0}; // @[AddRecFN.scala 73:58]
  wire [26:0] _close_alignedSigA_T_4 = 10'sh0 <= $signed(sDiffExps) & sDiffExps[0] ? _close_alignedSigA_T_3 : 27'h0; // @[AddRecFN.scala 73:12]
  wire [25:0] _close_alignedSigA_T_9 = {io_a_sig, 1'h0}; // @[AddRecFN.scala 74:58]
  wire [25:0] _close_alignedSigA_T_10 = _close_alignedSigA_T & ~sDiffExps[0] ? _close_alignedSigA_T_9 : 26'h0; // @[AddRecFN.scala 74:12]
  wire [26:0] _GEN_0 = {{1'd0}, _close_alignedSigA_T_10}; // @[AddRecFN.scala 73:68]
  wire [26:0] _close_alignedSigA_T_11 = _close_alignedSigA_T_4 | _GEN_0; // @[AddRecFN.scala 73:68]
  wire [24:0] _close_alignedSigA_T_13 = _modNatAlignDist_T ? io_a_sig : 25'h0; // @[AddRecFN.scala 75:12]
  wire [26:0] _GEN_1 = {{2'd0}, _close_alignedSigA_T_13}; // @[AddRecFN.scala 74:68]
  wire [26:0] _close_sSigSum_T = _close_alignedSigA_T_11 | _GEN_1; // @[AddRecFN.scala 76:43]
  wire [25:0] _close_sSigSum_T_2 = {io_b_sig, 1'h0}; // @[AddRecFN.scala 76:66]
  wire [26:0] _GEN_2 = {{1{_close_sSigSum_T_2[25]}},_close_sSigSum_T_2}; // @[AddRecFN.scala 76:50]
  wire [26:0] close_sSigSum = $signed(_close_sSigSum_T) - $signed(_GEN_2); // @[AddRecFN.scala 76:50]
  wire  _close_sigSum_T = $signed(close_sSigSum) < 27'sh0; // @[AddRecFN.scala 77:42]
  wire [26:0] _close_sigSum_T_3 = 27'sh0 - $signed(close_sSigSum); // @[AddRecFN.scala 77:49]
  wire [26:0] _close_sigSum_T_4 = $signed(close_sSigSum) < 27'sh0 ? $signed(_close_sigSum_T_3) : $signed(close_sSigSum); // @[AddRecFN.scala 77:27]
  wire [25:0] close_sigSum = _close_sigSum_T_4[25:0]; // @[AddRecFN.scala 77:79]
  wire  close_reduced2SigSum_reducedVec_0 = |close_sigSum[1:0]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_1 = |close_sigSum[3:2]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_2 = |close_sigSum[5:4]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_3 = |close_sigSum[7:6]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_4 = |close_sigSum[9:8]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_5 = |close_sigSum[11:10]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_6 = |close_sigSum[13:12]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_7 = |close_sigSum[15:14]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_8 = |close_sigSum[17:16]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_9 = |close_sigSum[19:18]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_10 = |close_sigSum[21:20]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_11 = |close_sigSum[23:22]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_12 = |close_sigSum[25:24]; // @[primitives.scala 106:57]
  wire [5:0] close_reduced2SigSum_lo = {close_reduced2SigSum_reducedVec_5,close_reduced2SigSum_reducedVec_4,
    close_reduced2SigSum_reducedVec_3,close_reduced2SigSum_reducedVec_2,close_reduced2SigSum_reducedVec_1,
    close_reduced2SigSum_reducedVec_0}; // @[primitives.scala 107:20]
  wire [12:0] close_reduced2SigSum = {close_reduced2SigSum_reducedVec_12,close_reduced2SigSum_reducedVec_11,
    close_reduced2SigSum_reducedVec_10,close_reduced2SigSum_reducedVec_9,close_reduced2SigSum_reducedVec_8,
    close_reduced2SigSum_reducedVec_7,close_reduced2SigSum_reducedVec_6,close_reduced2SigSum_lo}; // @[primitives.scala 107:20]
  wire [3:0] _close_normDistReduced2_T_13 = close_reduced2SigSum[1] ? 4'hb : 4'hc; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_14 = close_reduced2SigSum[2] ? 4'ha : _close_normDistReduced2_T_13; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_15 = close_reduced2SigSum[3] ? 4'h9 : _close_normDistReduced2_T_14; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_16 = close_reduced2SigSum[4] ? 4'h8 : _close_normDistReduced2_T_15; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_17 = close_reduced2SigSum[5] ? 4'h7 : _close_normDistReduced2_T_16; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_18 = close_reduced2SigSum[6] ? 4'h6 : _close_normDistReduced2_T_17; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_19 = close_reduced2SigSum[7] ? 4'h5 : _close_normDistReduced2_T_18; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_20 = close_reduced2SigSum[8] ? 4'h4 : _close_normDistReduced2_T_19; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_21 = close_reduced2SigSum[9] ? 4'h3 : _close_normDistReduced2_T_20; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_22 = close_reduced2SigSum[10] ? 4'h2 : _close_normDistReduced2_T_21; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_23 = close_reduced2SigSum[11] ? 4'h1 : _close_normDistReduced2_T_22; // @[Mux.scala 47:70]
  wire [3:0] close_normDistReduced2 = close_reduced2SigSum[12] ? 4'h0 : _close_normDistReduced2_T_23; // @[Mux.scala 47:70]
  wire [4:0] close_nearNormDist = {close_normDistReduced2, 1'h0}; // @[AddRecFN.scala 81:53]
  wire [56:0] _GEN_7 = {{31'd0}, close_sigSum}; // @[AddRecFN.scala 82:38]
  wire [56:0] _close_sigOut_T = _GEN_7 << close_nearNormDist; // @[AddRecFN.scala 82:38]
  wire [57:0] _close_sigOut_T_1 = {_close_sigOut_T, 1'h0}; // @[AddRecFN.scala 82:59]
  wire [26:0] close_sigOut = _close_sigOut_T_1[26:0]; // @[AddRecFN.scala 82:63]
  wire  close_totalCancellation = ~(|close_sigOut[26:25]); // @[AddRecFN.scala 83:35]
  wire  close_notTotalCancellation_signOut = io_a_sign ^ _close_sigSum_T; // @[AddRecFN.scala 84:56]
  wire  far_signOut = _modNatAlignDist_T ? effSignB : io_a_sign; // @[AddRecFN.scala 87:26]
  wire [24:0] _far_sigLarger_T_1 = _modNatAlignDist_T ? io_b_sig : io_a_sig; // @[AddRecFN.scala 88:29]
  wire [23:0] far_sigLarger = _far_sigLarger_T_1[23:0]; // @[AddRecFN.scala 88:66]
  wire [24:0] _far_sigSmaller_T_1 = _modNatAlignDist_T ? io_a_sig : io_b_sig; // @[AddRecFN.scala 89:29]
  wire [23:0] far_sigSmaller = _far_sigSmaller_T_1[23:0]; // @[AddRecFN.scala 89:66]
  wire [28:0] _far_mainAlignedSigSmaller_T = {far_sigSmaller, 5'h0}; // @[AddRecFN.scala 90:52]
  wire [28:0] far_mainAlignedSigSmaller = _far_mainAlignedSigSmaller_T >> alignDist; // @[AddRecFN.scala 90:56]
  wire [25:0] _far_reduced4SigSmaller_T = {far_sigSmaller, 2'h0}; // @[AddRecFN.scala 91:60]
  wire  far_reduced4SigSmaller_reducedVec_0 = |_far_reduced4SigSmaller_T[3:0]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_1 = |_far_reduced4SigSmaller_T[7:4]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_2 = |_far_reduced4SigSmaller_T[11:8]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_3 = |_far_reduced4SigSmaller_T[15:12]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_4 = |_far_reduced4SigSmaller_T[19:16]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_5 = |_far_reduced4SigSmaller_T[23:20]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_6 = |_far_reduced4SigSmaller_T[25:24]; // @[primitives.scala 123:57]
  wire [6:0] far_reduced4SigSmaller = {far_reduced4SigSmaller_reducedVec_6,far_reduced4SigSmaller_reducedVec_5,
    far_reduced4SigSmaller_reducedVec_4,far_reduced4SigSmaller_reducedVec_3,far_reduced4SigSmaller_reducedVec_2,
    far_reduced4SigSmaller_reducedVec_1,far_reduced4SigSmaller_reducedVec_0}; // @[primitives.scala 124:20]
  wire [8:0] far_roundExtraMask_shift = 9'sh100 >>> alignDist[4:2]; // @[primitives.scala 76:56]
  wire [6:0] far_roundExtraMask = {far_roundExtraMask_shift[1],far_roundExtraMask_shift[2],far_roundExtraMask_shift[3],
    far_roundExtraMask_shift[4],far_roundExtraMask_shift[5],far_roundExtraMask_shift[6],far_roundExtraMask_shift[7]}; // @[Cat.scala 33:92]
  wire [6:0] _far_alignedSigSmaller_T_3 = far_reduced4SigSmaller & far_roundExtraMask; // @[AddRecFN.scala 95:76]
  wire  _far_alignedSigSmaller_T_5 = |far_mainAlignedSigSmaller[2:0] | |_far_alignedSigSmaller_T_3; // @[AddRecFN.scala 95:49]
  wire [26:0] far_alignedSigSmaller = {far_mainAlignedSigSmaller[28:3],_far_alignedSigSmaller_T_5}; // @[Cat.scala 33:92]
  wire [26:0] _far_negAlignedSigSmaller_T = ~far_alignedSigSmaller; // @[AddRecFN.scala 97:62]
  wire [27:0] _far_negAlignedSigSmaller_T_1 = {1'h1,_far_negAlignedSigSmaller_T}; // @[Cat.scala 33:92]
  wire [27:0] far_negAlignedSigSmaller = _closeSubMags_T ? _far_negAlignedSigSmaller_T_1 : {{1'd0},
    far_alignedSigSmaller}; // @[AddRecFN.scala 97:39]
  wire [26:0] _far_sigSum_T = {far_sigLarger, 3'h0}; // @[AddRecFN.scala 98:36]
  wire [27:0] _GEN_3 = {{1'd0}, _far_sigSum_T}; // @[AddRecFN.scala 98:41]
  wire [27:0] _far_sigSum_T_2 = _GEN_3 + far_negAlignedSigSmaller; // @[AddRecFN.scala 98:41]
  wire [27:0] _GEN_4 = {{27'd0}, _closeSubMags_T}; // @[AddRecFN.scala 98:68]
  wire [27:0] far_sigSum = _far_sigSum_T_2 + _GEN_4; // @[AddRecFN.scala 98:68]
  wire [26:0] _GEN_5 = {{26'd0}, far_sigSum[0]}; // @[AddRecFN.scala 99:67]
  wire [26:0] _far_sigOut_T_2 = far_sigSum[27:1] | _GEN_5; // @[AddRecFN.scala 99:67]
  wire [27:0] _far_sigOut_T_3 = _closeSubMags_T ? far_sigSum : {{1'd0}, _far_sigOut_T_2}; // @[AddRecFN.scala 99:25]
  wire [26:0] far_sigOut = _far_sigOut_T_3[26:0]; // @[AddRecFN.scala 99:83]
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isInf & _closeSubMags_T; // @[AddRecFN.scala 102:57]
  wire  notNaN_isInfOut = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  wire  addZeros = io_a_isZero & io_b_isZero; // @[AddRecFN.scala 104:32]
  wire  notNaN_specialCase = notNaN_isInfOut | addZeros; // @[AddRecFN.scala 105:46]
  wire  _notNaN_signOut_T_1 = io_a_isInf & io_a_sign; // @[AddRecFN.scala 109:39]
  wire  _notNaN_signOut_T_2 = eqSigns & io_a_sign | _notNaN_signOut_T_1; // @[AddRecFN.scala 108:63]
  wire  _notNaN_signOut_T_3 = io_b_isInf & effSignB; // @[AddRecFN.scala 110:39]
  wire  _notNaN_signOut_T_4 = _notNaN_signOut_T_2 | _notNaN_signOut_T_3; // @[AddRecFN.scala 109:63]
  wire  _notNaN_signOut_T_9 = ~notNaN_specialCase; // @[AddRecFN.scala 112:10]
  wire  _notNaN_signOut_T_12 = ~notNaN_specialCase & closeSubMags & ~close_totalCancellation; // @[AddRecFN.scala 112:46]
  wire  _notNaN_signOut_T_13 = _notNaN_signOut_T_12 & close_notTotalCancellation_signOut; // @[AddRecFN.scala 113:38]
  wire  _notNaN_signOut_T_14 = _notNaN_signOut_T_4 | _notNaN_signOut_T_13; // @[AddRecFN.scala 111:63]
  wire  _notNaN_signOut_T_18 = _notNaN_signOut_T_9 & ~closeSubMags & far_signOut; // @[AddRecFN.scala 114:47]
  wire [9:0] _common_sExpOut_T_2 = closeSubMags | _modNatAlignDist_T ? $signed(io_b_sExp) : $signed(io_a_sExp); // @[AddRecFN.scala 116:13]
  wire [4:0] _common_sExpOut_T_3 = closeSubMags ? close_nearNormDist : {{4'd0}, _closeSubMags_T}; // @[AddRecFN.scala 117:18]
  wire [5:0] _common_sExpOut_T_4 = {1'b0,$signed(_common_sExpOut_T_3)}; // @[AddRecFN.scala 117:66]
  wire [9:0] _GEN_6 = {{4{_common_sExpOut_T_4[5]}},_common_sExpOut_T_4}; // @[AddRecFN.scala 117:13]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[AddRecFN.scala 121:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[AddRecFN.scala 125:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  assign io_rawOut_isZero = addZeros | ~notNaN_isInfOut & closeSubMags & close_totalCancellation; // @[AddRecFN.scala 106:37]
  assign io_rawOut_sign = _notNaN_signOut_T_14 | _notNaN_signOut_T_18; // @[AddRecFN.scala 113:77]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - $signed(_GEN_6); // @[AddRecFN.scala 117:13]
  assign io_rawOut_sig = closeSubMags ? close_sigOut : far_sigOut; // @[AddRecFN.scala 118:28]
endmodule
module AddRecFN(
  input         io_subOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  output [32:0] io_out
);
  wire  addRawFN__io_subOp; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_a_sExp; // @[AddRecFN.scala 147:26]
  wire [24:0] addRawFN__io_a_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_b_sExp; // @[AddRecFN.scala 147:26]
  wire [24:0] addRawFN__io_b_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_invalidExc; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 147:26]
  wire [26:0] addRawFN__io_rawOut_sig; // @[AddRecFN.scala 147:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[AddRecFN.scala 157:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[AddRecFN.scala 157:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[AddRecFN.scala 157:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[AddRecFN.scala 157:15]
  wire [8:0] addRawFN_io_a_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  addRawFN_io_a_isZero = addRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  addRawFN_io_a_isSpecial = addRawFN_io_a_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _addRawFN_io_a_out_sig_T = ~addRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _addRawFN_io_a_out_sig_T_1 = {1'h0,_addRawFN_io_a_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  wire [8:0] addRawFN_io_b_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  addRawFN_io_b_isZero = addRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  addRawFN_io_b_isSpecial = addRawFN_io_b_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _addRawFN_io_b_out_sig_T = ~addRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _addRawFN_io_b_out_sig_T_1 = {1'h0,_addRawFN_io_b_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  AddRawFN addRawFN_ ( // @[AddRecFN.scala 147:26]
    .io_subOp(addRawFN__io_subOp),
    .io_a_isNaN(addRawFN__io_a_isNaN),
    .io_a_isInf(addRawFN__io_a_isInf),
    .io_a_isZero(addRawFN__io_a_isZero),
    .io_a_sign(addRawFN__io_a_sign),
    .io_a_sExp(addRawFN__io_a_sExp),
    .io_a_sig(addRawFN__io_a_sig),
    .io_b_isNaN(addRawFN__io_b_isNaN),
    .io_b_isInf(addRawFN__io_b_isInf),
    .io_b_isZero(addRawFN__io_b_isZero),
    .io_b_sign(addRawFN__io_b_sign),
    .io_b_sExp(addRawFN__io_b_sExp),
    .io_b_sig(addRawFN__io_b_sig),
    .io_invalidExc(addRawFN__io_invalidExc),
    .io_rawOut_isNaN(addRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(addRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(addRawFN__io_rawOut_isZero),
    .io_rawOut_sign(addRawFN__io_rawOut_sign),
    .io_rawOut_sExp(addRawFN__io_rawOut_sExp),
    .io_rawOut_sig(addRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN_e8_s24 roundRawFNToRecFN ( // @[AddRecFN.scala 157:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[AddRecFN.scala 163:23]
  assign addRawFN__io_subOp = io_subOp; // @[AddRecFN.scala 149:30]
  assign addRawFN__io_a_isNaN = addRawFN_io_a_isSpecial & addRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_a_isInf = addRawFN_io_a_isSpecial & ~addRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign addRawFN__io_a_isZero = addRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign addRawFN__io_a_sign = io_a[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign addRawFN__io_a_sExp = {1'b0,$signed(addRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign addRawFN__io_a_sig = {_addRawFN_io_a_out_sig_T_1,io_a[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign addRawFN__io_b_isNaN = addRawFN_io_b_isSpecial & addRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_b_isInf = addRawFN_io_b_isSpecial & ~addRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign addRawFN__io_b_isZero = addRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign addRawFN__io_b_sign = io_b[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign addRawFN__io_b_sExp = {1'b0,$signed(addRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign addRawFN__io_b_sig = {_addRawFN_io_b_out_sig_T_1,io_b[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign roundRawFNToRecFN_io_invalidExc = addRawFN__io_invalidExc; // @[AddRecFN.scala 158:39]
  assign roundRawFNToRecFN_io_in_isNaN = addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isInf = addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isZero = addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sign = addRawFN__io_rawOut_sign; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sExp = addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sig = addRawFN__io_rawOut_sig; // @[AddRecFN.scala 160:39]
endmodule
module FP32Sub(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire  adder_io_subOp; // @[FPU.scala 45:23]
  wire [32:0] adder_io_a; // @[FPU.scala 45:23]
  wire [32:0] adder_io_b; // @[FPU.scala 45:23]
  wire [32:0] adder_io_out; // @[FPU.scala 45:23]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = adder_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = adder_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,adder_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  AddRecFN adder ( // @[FPU.scala 45:23]
    .io_subOp(adder_io_subOp),
    .io_a(adder_io_a),
    .io_b(adder_io_b),
    .io_out(adder_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign adder_io_subOp = 1'h1; // @[FPU.scala 52:20]
  assign adder_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign adder_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module FP32radianCaclulator(
  input         clock,
  input         reset,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_m,
  input  [31:0] io_baseIndex,
  input  [31:0] io_TwoDivD,
  output [31:0] io_out,
  output        io_ENout,
  output [31:0] io_xFWD_0,
  output [31:0] io_xFWD_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] Int64ToFP32_io_inInt; // @[RoPEModuleFP32.scala 36:29]
  wire [31:0] Int64ToFP32_io_outIEEE; // @[RoPEModuleFP32.scala 36:29]
  wire [31:0] FP32Mult0_io_a; // @[RoPEModuleFP32.scala 41:27]
  wire [31:0] FP32Mult0_io_b; // @[RoPEModuleFP32.scala 41:27]
  wire [31:0] FP32Mult0_io_result; // @[RoPEModuleFP32.scala 41:27]
  wire [31:0] FP32DivPOW2_io_a; // @[RoPEModuleFP32.scala 47:29]
  wire [31:0] FP32DivPOW2_io_result; // @[RoPEModuleFP32.scala 47:29]
  wire [31:0] FP32Mult1_io_a; // @[RoPEModuleFP32.scala 54:27]
  wire [31:0] FP32Mult1_io_b; // @[RoPEModuleFP32.scala 54:27]
  wire [31:0] FP32Mult1_io_result; // @[RoPEModuleFP32.scala 54:27]
  wire [31:0] FP32Sub_io_a; // @[RoPEModuleFP32.scala 64:25]
  wire [31:0] FP32Sub_io_b; // @[RoPEModuleFP32.scala 64:25]
  wire [31:0] FP32Sub_io_result; // @[RoPEModuleFP32.scala 64:25]
  wire [32:0] _stage1Reg_T = {{1'd0}, io_baseIndex}; // @[RoPEModuleFP32.scala 17:89]
  reg [63:0] stage1Reg_0; // @[RoPEModuleFP32.scala 17:28]
  reg [63:0] stage1Reg_1; // @[RoPEModuleFP32.scala 17:28]
  reg [63:0] stage1Reg_2; // @[RoPEModuleFP32.scala 17:28]
  reg [63:0] stage1Reg_3; // @[RoPEModuleFP32.scala 17:28]
  reg [31:0] stage2Reg_0; // @[RoPEModuleFP32.scala 19:28]
  reg [31:0] stage2Reg_1; // @[RoPEModuleFP32.scala 19:28]
  reg [31:0] stage2Reg_2; // @[RoPEModuleFP32.scala 19:28]
  reg [31:0] stage2Reg_3; // @[RoPEModuleFP32.scala 19:28]
  reg [31:0] stage3Reg_0; // @[RoPEModuleFP32.scala 20:28]
  reg [31:0] stage3Reg_1; // @[RoPEModuleFP32.scala 20:28]
  reg [31:0] stage3Reg_2; // @[RoPEModuleFP32.scala 20:28]
  reg [31:0] stage4Reg_0; // @[RoPEModuleFP32.scala 21:28]
  reg [31:0] stage4Reg_1; // @[RoPEModuleFP32.scala 21:28]
  reg [31:0] stage4Reg_2; // @[RoPEModuleFP32.scala 21:28]
  reg [31:0] stage5Reg_0; // @[RoPEModuleFP32.scala 22:28]
  reg [31:0] stage5Reg_1; // @[RoPEModuleFP32.scala 22:28]
  reg [31:0] stage5Reg_2; // @[RoPEModuleFP32.scala 22:28]
  reg [31:0] stage5Reg_3; // @[RoPEModuleFP32.scala 22:28]
  reg [31:0] stage6Reg_0; // @[RoPEModuleFP32.scala 23:28]
  reg [31:0] stage6Reg_1; // @[RoPEModuleFP32.scala 23:28]
  reg [31:0] stage6Reg_2; // @[RoPEModuleFP32.scala 23:28]
  reg  enReg_0; // @[RoPEModuleFP32.scala 24:24]
  reg  enReg_1; // @[RoPEModuleFP32.scala 24:24]
  reg  enReg_2; // @[RoPEModuleFP32.scala 24:24]
  reg  enReg_3; // @[RoPEModuleFP32.scala 24:24]
  reg  enReg_4; // @[RoPEModuleFP32.scala 24:24]
  reg  enReg_5; // @[RoPEModuleFP32.scala 24:24]
  reg [31:0] delayedMThetaI; // @[RoPEModuleFP32.scala 60:33]
  wire [63:0] _WIRE__3 = {{32'd0}, Int64ToFP32_io_outIEEE}; // @[RoPEModuleFP32.scala 38:{25,25}]
  wire [31:0] _WIRE_1_2 = FP32Mult0_io_result; // @[RoPEModuleFP32.scala 44:{25,25}]
  wire [31:0] _WIRE_2_2 = FP32DivPOW2_io_result; // @[RoPEModuleFP32.scala 51:{25,25}]
  wire [31:0] _WIRE_3_3 = FP32Mult1_io_result; // @[RoPEModuleFP32.scala 57:{25,25}]
  wire [31:0] _WIRE_4_2 = FP32Sub_io_result; // @[RoPEModuleFP32.scala 68:{25,25}]
  wire [63:0] _GEN_0 = reset ? 64'h0 : stage1Reg_0; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
  wire [63:0] _GEN_1 = reset ? 64'h0 : stage1Reg_1; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
  wire [63:0] _GEN_2 = reset ? 64'h0 : stage1Reg_2; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
  wire [63:0] _GEN_3 = reset ? 64'h0 : _WIRE__3; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
  Int64ToFP32 Int64ToFP32 ( // @[RoPEModuleFP32.scala 36:29]
    .io_inInt(Int64ToFP32_io_inInt),
    .io_outIEEE(Int64ToFP32_io_outIEEE)
  );
  FP32Multiplier FP32Mult0 ( // @[RoPEModuleFP32.scala 41:27]
    .io_a(FP32Mult0_io_a),
    .io_b(FP32Mult0_io_b),
    .io_result(FP32Mult0_io_result)
  );
  FP32DivPOW2INT FP32DivPOW2 ( // @[RoPEModuleFP32.scala 47:29]
    .io_a(FP32DivPOW2_io_a),
    .io_result(FP32DivPOW2_io_result)
  );
  FP32Multiplier FP32Mult1 ( // @[RoPEModuleFP32.scala 54:27]
    .io_a(FP32Mult1_io_a),
    .io_b(FP32Mult1_io_b),
    .io_result(FP32Mult1_io_result)
  );
  FP32Sub FP32Sub ( // @[RoPEModuleFP32.scala 64:25]
    .io_a(FP32Sub_io_a),
    .io_b(FP32Sub_io_b),
    .io_result(FP32Sub_io_result)
  );
  assign io_out = enReg_5 ? stage6Reg_2 : 32'h0; // @[RoPEModuleFP32.scala 71:22]
  assign io_ENout = enReg_5; // @[RoPEModuleFP32.scala 74:16]
  assign io_xFWD_0 = enReg_5 ? stage6Reg_0 : 32'h0; // @[RoPEModuleFP32.scala 72:22]
  assign io_xFWD_1 = enReg_5 ? stage6Reg_1 : 32'h0; // @[RoPEModuleFP32.scala 73:22]
  assign Int64ToFP32_io_inInt = stage1Reg_3; // @[RoPEModuleFP32.scala 37:42]
  assign FP32Mult0_io_a = stage2Reg_3; // @[RoPEModuleFP32.scala 42:20]
  assign FP32Mult0_io_b = stage2Reg_2; // @[RoPEModuleFP32.scala 43:20]
  assign FP32DivPOW2_io_a = stage3Reg_2; // @[RoPEModuleFP32.scala 48:22]
  assign FP32Mult1_io_a = stage4Reg_2; // @[RoPEModuleFP32.scala 55:20]
  assign FP32Mult1_io_b = 32'h40000000; // @[RoPEModuleFP32.scala 56:20]
  assign FP32Sub_io_a = delayedMThetaI; // @[RoPEModuleFP32.scala 66:18]
  assign FP32Sub_io_b = stage5Reg_3; // @[RoPEModuleFP32.scala 67:18]
  always @(posedge clock) begin
    stage1Reg_0 <= {{32'd0}, io_x_0}; // @[RoPEModuleFP32.scala 17:{36,36}]
    stage1Reg_1 <= {{32'd0}, io_x_1}; // @[RoPEModuleFP32.scala 17:{36,36}]
    stage1Reg_2 <= {{32'd0}, io_TwoDivD}; // @[RoPEModuleFP32.scala 17:{36,36}]
    stage1Reg_3 <= io_m * _stage1Reg_T[31:0]; // @[RoPEModuleFP32.scala 17:73]
    stage2Reg_0 <= _GEN_0[31:0]; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
    stage2Reg_1 <= _GEN_1[31:0]; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
    stage2Reg_2 <= _GEN_2[31:0]; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
    stage2Reg_3 <= _GEN_3[31:0]; // @[RoPEModuleFP32.scala 19:{28,28} 38:15]
    if (reset) begin // @[RoPEModuleFP32.scala 20:28]
      stage3Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 20:28]
    end else begin
      stage3Reg_0 <= stage2Reg_0; // @[RoPEModuleFP32.scala 44:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 20:28]
      stage3Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 20:28]
    end else begin
      stage3Reg_1 <= stage2Reg_1; // @[RoPEModuleFP32.scala 44:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 20:28]
      stage3Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 20:28]
    end else begin
      stage3Reg_2 <= _WIRE_1_2; // @[RoPEModuleFP32.scala 44:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 21:28]
      stage4Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 21:28]
    end else begin
      stage4Reg_0 <= stage3Reg_0; // @[RoPEModuleFP32.scala 51:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 21:28]
      stage4Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 21:28]
    end else begin
      stage4Reg_1 <= stage3Reg_1; // @[RoPEModuleFP32.scala 51:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 21:28]
      stage4Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 21:28]
    end else begin
      stage4Reg_2 <= _WIRE_2_2; // @[RoPEModuleFP32.scala 51:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 22:28]
      stage5Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 22:28]
    end else begin
      stage5Reg_0 <= stage4Reg_0; // @[RoPEModuleFP32.scala 57:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 22:28]
      stage5Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 22:28]
    end else begin
      stage5Reg_1 <= stage4Reg_1; // @[RoPEModuleFP32.scala 57:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 22:28]
      stage5Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 22:28]
    end else begin
      stage5Reg_2 <= stage3Reg_2; // @[RoPEModuleFP32.scala 57:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 22:28]
      stage5Reg_3 <= 32'h0; // @[RoPEModuleFP32.scala 22:28]
    end else begin
      stage5Reg_3 <= _WIRE_3_3; // @[RoPEModuleFP32.scala 57:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 23:28]
      stage6Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 23:28]
    end else begin
      stage6Reg_0 <= stage5Reg_0; // @[RoPEModuleFP32.scala 68:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 23:28]
      stage6Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 23:28]
    end else begin
      stage6Reg_1 <= stage5Reg_1; // @[RoPEModuleFP32.scala 68:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 23:28]
      stage6Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 23:28]
    end else begin
      stage6Reg_2 <= _WIRE_4_2; // @[RoPEModuleFP32.scala 68:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_0 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_0 <= io_EN; // @[RoPEModuleFP32.scala 27:14]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_1 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_1 <= enReg_0; // @[RoPEModuleFP32.scala 29:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_2 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_2 <= enReg_1; // @[RoPEModuleFP32.scala 29:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_3 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_3 <= enReg_2; // @[RoPEModuleFP32.scala 29:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_4 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_4 <= enReg_3; // @[RoPEModuleFP32.scala 29:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 24:24]
      enReg_5 <= 1'h0; // @[RoPEModuleFP32.scala 24:24]
    end else begin
      enReg_5 <= enReg_4; // @[RoPEModuleFP32.scala 29:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 60:33]
      delayedMThetaI <= 32'h0; // @[RoPEModuleFP32.scala 60:33]
    end else begin
      delayedMThetaI <= stage5Reg_2; // @[RoPEModuleFP32.scala 61:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  stage1Reg_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  stage1Reg_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  stage1Reg_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  stage1Reg_3 = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  stage2Reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stage2Reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stage2Reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage2Reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage3Reg_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage3Reg_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stage3Reg_2 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stage4Reg_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stage4Reg_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  stage4Reg_2 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stage5Reg_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stage5Reg_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  stage5Reg_2 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  stage5Reg_3 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  stage6Reg_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  stage6Reg_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stage6Reg_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  enReg_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  enReg_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  enReg_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  enReg_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  enReg_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  enReg_5 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  delayedMThetaI = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP32toINT32(
  input  [31:0] io_ieee754,
  output [31:0] io_int32
);
  wire  sign = io_ieee754[31]; // @[FPU.scala 242:24]
  wire [7:0] exponent = io_ieee754[30:23]; // @[FPU.scala 243:37]
  wire [22:0] mantissa = io_ieee754[22:0]; // @[FPU.scala 244:28]
  wire [23:0] mantissaWithLeadingOne = {1'h1,mantissa}; // @[Cat.scala 33:92]
  wire [7:0] trueExponent = $signed(exponent) - 8'sh7f; // @[FPU.scala 250:31]
  wire [7:0] shiftAmount = $signed(trueExponent) - 8'sh17; // @[FPU.scala 253:34]
  wire [7:0] _shiftedMantissa_T_1 = $signed(trueExponent) - 8'sh17; // @[FPU.scala 257:43]
  wire [278:0] _GEN_1 = {{255'd0}, mantissaWithLeadingOne}; // @[FPU.scala 257:28]
  wire [278:0] _shiftedMantissa_T_2 = _GEN_1 << _shiftedMantissa_T_1; // @[FPU.scala 257:28]
  wire [7:0] _shiftedMantissa_T_5 = 8'h0 - _shiftedMantissa_T_1; // @[FPU.scala 258:31]
  wire [23:0] _shiftedMantissa_T_6 = mantissaWithLeadingOne >> _shiftedMantissa_T_5; // @[FPU.scala 258:28]
  wire [278:0] _result_T_1 = $signed(shiftAmount) >= 8'sh0 ? _shiftedMantissa_T_2 : {{255'd0}, _shiftedMantissa_T_6}; // @[FPU.scala 261:50]
  wire [278:0] _result_T_5 = 279'sh0 - $signed(_result_T_1); // @[FPU.scala 261:58]
  wire [278:0] result = ~sign ? $signed(_result_T_1) : $signed(_result_T_5); // @[FPU.scala 261:19]
  assign io_int32 = result[31:0]; // @[FPU.scala 264:12]
endmodule
module IndexCalculator(
  input         io_EN,
  input  [31:0] io_angle,
  output [31:0] io_cosIndex,
  output [31:0] io_sinIndex,
  output        io_cosSign,
  output        io_sinSign,
  output        io_ENout
);
  wire [31:0] FP32Mult_io_a; // @[sincosLUT.scala 18:32]
  wire [31:0] FP32Mult_io_b; // @[sincosLUT.scala 18:32]
  wire [31:0] FP32Mult_io_result; // @[sincosLUT.scala 18:32]
  wire [31:0] FP32Truncate_io_in; // @[sincosLUT.scala 19:32]
  wire [31:0] FP32Truncate_io_out; // @[sincosLUT.scala 19:32]
  wire [31:0] FP32toINT32_io_ieee754; // @[sincosLUT.scala 20:32]
  wire [31:0] FP32toINT32_io_int32; // @[sincosLUT.scala 20:32]
  wire [31:0] _cosIndexWire_T_1 = 32'h800 - FP32toINT32_io_int32; // @[sincosLUT.scala 55:28]
  wire  _T_2 = FP32toINT32_io_int32 <= 32'hc00; // @[sincosLUT.scala 59:22]
  wire [31:0] _cosIndexWire_T_3 = FP32toINT32_io_int32 - 32'h800; // @[sincosLUT.scala 60:31]
  wire [31:0] _cosIndexWire_T_5 = 32'h1000 - FP32toINT32_io_int32; // @[sincosLUT.scala 65:34]
  wire [31:0] _GEN_0 = FP32toINT32_io_int32 <= 32'hc00 ? _cosIndexWire_T_3 : _cosIndexWire_T_5; // @[sincosLUT.scala 59:39 60:22 65:22]
  wire [31:0] _GEN_4 = FP32toINT32_io_int32 <= 32'h800 ? _cosIndexWire_T_1 : _GEN_0; // @[sincosLUT.scala 54:29 55:22]
  wire  _GEN_6 = FP32toINT32_io_int32 <= 32'h800 | _T_2; // @[sincosLUT.scala 54:29 57:22]
  wire  _GEN_7 = FP32toINT32_io_int32 <= 32'h800 ? 1'h0 : 1'h1; // @[sincosLUT.scala 54:29 58:22]
  wire [31:0] cosIndexWire = FP32toINT32_io_int32 <= 32'h400 ? FP32toINT32_io_int32 : _GEN_4; // @[sincosLUT.scala 49:27 50:22]
  wire  cosSignWire = FP32toINT32_io_int32 <= 32'h400 ? 1'h0 : _GEN_6; // @[sincosLUT.scala 49:27 52:22]
  wire  sinSignWire = FP32toINT32_io_int32 <= 32'h400 ? 1'h0 : _GEN_7; // @[sincosLUT.scala 49:27 53:22]
  FP32Multiplier FP32Mult ( // @[sincosLUT.scala 18:32]
    .io_a(FP32Mult_io_a),
    .io_b(FP32Mult_io_b),
    .io_result(FP32Mult_io_result)
  );
  FP32Truncate FP32Truncate ( // @[sincosLUT.scala 19:32]
    .io_in(FP32Truncate_io_in),
    .io_out(FP32Truncate_io_out)
  );
  FP32toINT32 FP32toINT32 ( // @[sincosLUT.scala 20:32]
    .io_ieee754(FP32toINT32_io_ieee754),
    .io_int32(FP32toINT32_io_int32)
  );
  assign io_cosIndex = io_EN ? cosIndexWire : 32'h0; // @[sincosLUT.scala 72:23]
  assign io_sinIndex = io_EN ? cosIndexWire : 32'h0; // @[sincosLUT.scala 73:23]
  assign io_cosSign = io_EN & cosSignWire; // @[sincosLUT.scala 74:23]
  assign io_sinSign = io_EN & sinSignWire; // @[sincosLUT.scala 75:23]
  assign io_ENout = io_EN; // @[sincosLUT.scala 76:17]
  assign FP32Mult_io_a = io_angle; // @[sincosLUT.scala 22:19]
  assign FP32Mult_io_b = 32'h45000000; // @[sincosLUT.scala 23:19]
  assign FP32Truncate_io_in = FP32Mult_io_result; // @[sincosLUT.scala 26:24]
  assign FP32toINT32_io_ieee754 = FP32Truncate_io_out; // @[sincosLUT.scala 29:28]
endmodule
module CosLUT(
  input         io_EN,
  input  [31:0] io_cosIndex,
  input  [31:0] io_sinIndex,
  output [31:0] io_sinOut,
  output [31:0] io_cosOut,
  output        io_ENout
);
  wire [29:0] _GEN_1 = 11'h1 == io_cosIndex[10:0] ? 30'h3f7fffec : 30'h3f800000; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_2 = 11'h2 == io_cosIndex[10:0] ? 30'h3f7fffb1 : _GEN_1; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_3 = 11'h3 == io_cosIndex[10:0] ? 30'h3f7fff4e : _GEN_2; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_4 = 11'h4 == io_cosIndex[10:0] ? 30'h3f7ffec4 : _GEN_3; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_5 = 11'h5 == io_cosIndex[10:0] ? 30'h3f7ffe12 : _GEN_4; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_6 = 11'h6 == io_cosIndex[10:0] ? 30'h3f7ffd39 : _GEN_5; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_7 = 11'h7 == io_cosIndex[10:0] ? 30'h3f7ffc38 : _GEN_6; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_8 = 11'h8 == io_cosIndex[10:0] ? 30'h3f7ffb10 : _GEN_7; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_9 = 11'h9 == io_cosIndex[10:0] ? 30'h3f7ff9c0 : _GEN_8; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_10 = 11'ha == io_cosIndex[10:0] ? 30'h3f7ff849 : _GEN_9; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_11 = 11'hb == io_cosIndex[10:0] ? 30'h3f7ff6aa : _GEN_10; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_12 = 11'hc == io_cosIndex[10:0] ? 30'h3f7ff4e4 : _GEN_11; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_13 = 11'hd == io_cosIndex[10:0] ? 30'h3f7ff2f7 : _GEN_12; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_14 = 11'he == io_cosIndex[10:0] ? 30'h3f7ff0e1 : _GEN_13; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_15 = 11'hf == io_cosIndex[10:0] ? 30'h3f7feea5 : _GEN_14; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_16 = 11'h10 == io_cosIndex[10:0] ? 30'h3f7fec41 : _GEN_15; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_17 = 11'h11 == io_cosIndex[10:0] ? 30'h3f7fe9b5 : _GEN_16; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_18 = 11'h12 == io_cosIndex[10:0] ? 30'h3f7fe702 : _GEN_17; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_19 = 11'h13 == io_cosIndex[10:0] ? 30'h3f7fe427 : _GEN_18; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_20 = 11'h14 == io_cosIndex[10:0] ? 30'h3f7fe125 : _GEN_19; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_21 = 11'h15 == io_cosIndex[10:0] ? 30'h3f7fddfc : _GEN_20; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_22 = 11'h16 == io_cosIndex[10:0] ? 30'h3f7fdaaa : _GEN_21; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_23 = 11'h17 == io_cosIndex[10:0] ? 30'h3f7fd732 : _GEN_22; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_24 = 11'h18 == io_cosIndex[10:0] ? 30'h3f7fd392 : _GEN_23; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_25 = 11'h19 == io_cosIndex[10:0] ? 30'h3f7fcfca : _GEN_24; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_26 = 11'h1a == io_cosIndex[10:0] ? 30'h3f7fcbdc : _GEN_25; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_27 = 11'h1b == io_cosIndex[10:0] ? 30'h3f7fc7c5 : _GEN_26; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_28 = 11'h1c == io_cosIndex[10:0] ? 30'h3f7fc387 : _GEN_27; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_29 = 11'h1d == io_cosIndex[10:0] ? 30'h3f7fbf22 : _GEN_28; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_30 = 11'h1e == io_cosIndex[10:0] ? 30'h3f7fba95 : _GEN_29; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_31 = 11'h1f == io_cosIndex[10:0] ? 30'h3f7fb5e1 : _GEN_30; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_32 = 11'h20 == io_cosIndex[10:0] ? 30'h3f7fb105 : _GEN_31; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_33 = 11'h21 == io_cosIndex[10:0] ? 30'h3f7fac02 : _GEN_32; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_34 = 11'h22 == io_cosIndex[10:0] ? 30'h3f7fa6d8 : _GEN_33; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_35 = 11'h23 == io_cosIndex[10:0] ? 30'h3f7fa185 : _GEN_34; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_36 = 11'h24 == io_cosIndex[10:0] ? 30'h3f7f9c0c : _GEN_35; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_37 = 11'h25 == io_cosIndex[10:0] ? 30'h3f7f966b : _GEN_36; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_38 = 11'h26 == io_cosIndex[10:0] ? 30'h3f7f90a3 : _GEN_37; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_39 = 11'h27 == io_cosIndex[10:0] ? 30'h3f7f8ab3 : _GEN_38; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_40 = 11'h28 == io_cosIndex[10:0] ? 30'h3f7f849c : _GEN_39; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_41 = 11'h29 == io_cosIndex[10:0] ? 30'h3f7f7e5d : _GEN_40; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_42 = 11'h2a == io_cosIndex[10:0] ? 30'h3f7f77f7 : _GEN_41; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_43 = 11'h2b == io_cosIndex[10:0] ? 30'h3f7f716a : _GEN_42; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_44 = 11'h2c == io_cosIndex[10:0] ? 30'h3f7f6ab5 : _GEN_43; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_45 = 11'h2d == io_cosIndex[10:0] ? 30'h3f7f63d8 : _GEN_44; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_46 = 11'h2e == io_cosIndex[10:0] ? 30'h3f7f5cd5 : _GEN_45; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_47 = 11'h2f == io_cosIndex[10:0] ? 30'h3f7f55aa : _GEN_46; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_48 = 11'h30 == io_cosIndex[10:0] ? 30'h3f7f4e57 : _GEN_47; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_49 = 11'h31 == io_cosIndex[10:0] ? 30'h3f7f46dd : _GEN_48; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_50 = 11'h32 == io_cosIndex[10:0] ? 30'h3f7f3f3c : _GEN_49; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_51 = 11'h33 == io_cosIndex[10:0] ? 30'h3f7f3773 : _GEN_50; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_52 = 11'h34 == io_cosIndex[10:0] ? 30'h3f7f2f83 : _GEN_51; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_53 = 11'h35 == io_cosIndex[10:0] ? 30'h3f7f276c : _GEN_52; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_54 = 11'h36 == io_cosIndex[10:0] ? 30'h3f7f1f2d : _GEN_53; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_55 = 11'h37 == io_cosIndex[10:0] ? 30'h3f7f16c7 : _GEN_54; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_56 = 11'h38 == io_cosIndex[10:0] ? 30'h3f7f0e3a : _GEN_55; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_57 = 11'h39 == io_cosIndex[10:0] ? 30'h3f7f0585 : _GEN_56; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_58 = 11'h3a == io_cosIndex[10:0] ? 30'h3f7efca9 : _GEN_57; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_59 = 11'h3b == io_cosIndex[10:0] ? 30'h3f7ef3a5 : _GEN_58; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_60 = 11'h3c == io_cosIndex[10:0] ? 30'h3f7eea7a : _GEN_59; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_61 = 11'h3d == io_cosIndex[10:0] ? 30'h3f7ee128 : _GEN_60; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_62 = 11'h3e == io_cosIndex[10:0] ? 30'h3f7ed7af : _GEN_61; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_63 = 11'h3f == io_cosIndex[10:0] ? 30'h3f7ece0e : _GEN_62; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_64 = 11'h40 == io_cosIndex[10:0] ? 30'h3f7ec446 : _GEN_63; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_65 = 11'h41 == io_cosIndex[10:0] ? 30'h3f7eba56 : _GEN_64; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_66 = 11'h42 == io_cosIndex[10:0] ? 30'h3f7eb03f : _GEN_65; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_67 = 11'h43 == io_cosIndex[10:0] ? 30'h3f7ea601 : _GEN_66; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_68 = 11'h44 == io_cosIndex[10:0] ? 30'h3f7e9b9c : _GEN_67; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_69 = 11'h45 == io_cosIndex[10:0] ? 30'h3f7e9110 : _GEN_68; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_70 = 11'h46 == io_cosIndex[10:0] ? 30'h3f7e865c : _GEN_69; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_71 = 11'h47 == io_cosIndex[10:0] ? 30'h3f7e7b80 : _GEN_70; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_72 = 11'h48 == io_cosIndex[10:0] ? 30'h3f7e707e : _GEN_71; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_73 = 11'h49 == io_cosIndex[10:0] ? 30'h3f7e6554 : _GEN_72; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_74 = 11'h4a == io_cosIndex[10:0] ? 30'h3f7e5a03 : _GEN_73; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_75 = 11'h4b == io_cosIndex[10:0] ? 30'h3f7e4e8b : _GEN_74; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_76 = 11'h4c == io_cosIndex[10:0] ? 30'h3f7e42ec : _GEN_75; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_77 = 11'h4d == io_cosIndex[10:0] ? 30'h3f7e3725 : _GEN_76; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_78 = 11'h4e == io_cosIndex[10:0] ? 30'h3f7e2b37 : _GEN_77; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_79 = 11'h4f == io_cosIndex[10:0] ? 30'h3f7e1f22 : _GEN_78; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_80 = 11'h50 == io_cosIndex[10:0] ? 30'h3f7e12e6 : _GEN_79; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_81 = 11'h51 == io_cosIndex[10:0] ? 30'h3f7e0682 : _GEN_80; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_82 = 11'h52 == io_cosIndex[10:0] ? 30'h3f7df9f8 : _GEN_81; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_83 = 11'h53 == io_cosIndex[10:0] ? 30'h3f7ded46 : _GEN_82; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_84 = 11'h54 == io_cosIndex[10:0] ? 30'h3f7de06d : _GEN_83; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_85 = 11'h55 == io_cosIndex[10:0] ? 30'h3f7dd36d : _GEN_84; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_86 = 11'h56 == io_cosIndex[10:0] ? 30'h3f7dc645 : _GEN_85; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_87 = 11'h57 == io_cosIndex[10:0] ? 30'h3f7db8f7 : _GEN_86; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_88 = 11'h58 == io_cosIndex[10:0] ? 30'h3f7dab81 : _GEN_87; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_89 = 11'h59 == io_cosIndex[10:0] ? 30'h3f7d9de4 : _GEN_88; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_90 = 11'h5a == io_cosIndex[10:0] ? 30'h3f7d9020 : _GEN_89; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_91 = 11'h5b == io_cosIndex[10:0] ? 30'h3f7d8235 : _GEN_90; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_92 = 11'h5c == io_cosIndex[10:0] ? 30'h3f7d7423 : _GEN_91; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_93 = 11'h5d == io_cosIndex[10:0] ? 30'h3f7d65ea : _GEN_92; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_94 = 11'h5e == io_cosIndex[10:0] ? 30'h3f7d5789 : _GEN_93; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_95 = 11'h5f == io_cosIndex[10:0] ? 30'h3f7d4902 : _GEN_94; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_96 = 11'h60 == io_cosIndex[10:0] ? 30'h3f7d3a53 : _GEN_95; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_97 = 11'h61 == io_cosIndex[10:0] ? 30'h3f7d2b7e : _GEN_96; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_98 = 11'h62 == io_cosIndex[10:0] ? 30'h3f7d1c81 : _GEN_97; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_99 = 11'h63 == io_cosIndex[10:0] ? 30'h3f7d0d5d : _GEN_98; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_100 = 11'h64 == io_cosIndex[10:0] ? 30'h3f7cfe13 : _GEN_99; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_101 = 11'h65 == io_cosIndex[10:0] ? 30'h3f7ceea1 : _GEN_100; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_102 = 11'h66 == io_cosIndex[10:0] ? 30'h3f7cdf08 : _GEN_101; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_103 = 11'h67 == io_cosIndex[10:0] ? 30'h3f7ccf48 : _GEN_102; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_104 = 11'h68 == io_cosIndex[10:0] ? 30'h3f7cbf61 : _GEN_103; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_105 = 11'h69 == io_cosIndex[10:0] ? 30'h3f7caf53 : _GEN_104; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_106 = 11'h6a == io_cosIndex[10:0] ? 30'h3f7c9f1f : _GEN_105; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_107 = 11'h6b == io_cosIndex[10:0] ? 30'h3f7c8ec3 : _GEN_106; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_108 = 11'h6c == io_cosIndex[10:0] ? 30'h3f7c7e40 : _GEN_107; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_109 = 11'h6d == io_cosIndex[10:0] ? 30'h3f7c6d96 : _GEN_108; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_110 = 11'h6e == io_cosIndex[10:0] ? 30'h3f7c5cc6 : _GEN_109; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_111 = 11'h6f == io_cosIndex[10:0] ? 30'h3f7c4bce : _GEN_110; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_112 = 11'h70 == io_cosIndex[10:0] ? 30'h3f7c3aaf : _GEN_111; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_113 = 11'h71 == io_cosIndex[10:0] ? 30'h3f7c296a : _GEN_112; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_114 = 11'h72 == io_cosIndex[10:0] ? 30'h3f7c17fe : _GEN_113; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_115 = 11'h73 == io_cosIndex[10:0] ? 30'h3f7c066a : _GEN_114; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_116 = 11'h74 == io_cosIndex[10:0] ? 30'h3f7bf4b0 : _GEN_115; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_117 = 11'h75 == io_cosIndex[10:0] ? 30'h3f7be2cf : _GEN_116; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_118 = 11'h76 == io_cosIndex[10:0] ? 30'h3f7bd0c7 : _GEN_117; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_119 = 11'h77 == io_cosIndex[10:0] ? 30'h3f7bbe99 : _GEN_118; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_120 = 11'h78 == io_cosIndex[10:0] ? 30'h3f7bac43 : _GEN_119; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_121 = 11'h79 == io_cosIndex[10:0] ? 30'h3f7b99c7 : _GEN_120; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_122 = 11'h7a == io_cosIndex[10:0] ? 30'h3f7b8723 : _GEN_121; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_123 = 11'h7b == io_cosIndex[10:0] ? 30'h3f7b7459 : _GEN_122; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_124 = 11'h7c == io_cosIndex[10:0] ? 30'h3f7b6169 : _GEN_123; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_125 = 11'h7d == io_cosIndex[10:0] ? 30'h3f7b4e51 : _GEN_124; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_126 = 11'h7e == io_cosIndex[10:0] ? 30'h3f7b3b13 : _GEN_125; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_127 = 11'h7f == io_cosIndex[10:0] ? 30'h3f7b27ad : _GEN_126; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_128 = 11'h80 == io_cosIndex[10:0] ? 30'h3f7b1422 : _GEN_127; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_129 = 11'h81 == io_cosIndex[10:0] ? 30'h3f7b006f : _GEN_128; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_130 = 11'h82 == io_cosIndex[10:0] ? 30'h3f7aec96 : _GEN_129; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_131 = 11'h83 == io_cosIndex[10:0] ? 30'h3f7ad895 : _GEN_130; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_132 = 11'h84 == io_cosIndex[10:0] ? 30'h3f7ac46f : _GEN_131; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_133 = 11'h85 == io_cosIndex[10:0] ? 30'h3f7ab021 : _GEN_132; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_134 = 11'h86 == io_cosIndex[10:0] ? 30'h3f7a9bad : _GEN_133; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_135 = 11'h87 == io_cosIndex[10:0] ? 30'h3f7a8712 : _GEN_134; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_136 = 11'h88 == io_cosIndex[10:0] ? 30'h3f7a7251 : _GEN_135; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_137 = 11'h89 == io_cosIndex[10:0] ? 30'h3f7a5d69 : _GEN_136; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_138 = 11'h8a == io_cosIndex[10:0] ? 30'h3f7a485a : _GEN_137; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_139 = 11'h8b == io_cosIndex[10:0] ? 30'h3f7a3325 : _GEN_138; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_140 = 11'h8c == io_cosIndex[10:0] ? 30'h3f7a1dc9 : _GEN_139; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_141 = 11'h8d == io_cosIndex[10:0] ? 30'h3f7a0846 : _GEN_140; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_142 = 11'h8e == io_cosIndex[10:0] ? 30'h3f79f29d : _GEN_141; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_143 = 11'h8f == io_cosIndex[10:0] ? 30'h3f79dccd : _GEN_142; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_144 = 11'h90 == io_cosIndex[10:0] ? 30'h3f79c6d7 : _GEN_143; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_145 = 11'h91 == io_cosIndex[10:0] ? 30'h3f79b0ba : _GEN_144; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_146 = 11'h92 == io_cosIndex[10:0] ? 30'h3f799a77 : _GEN_145; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_147 = 11'h93 == io_cosIndex[10:0] ? 30'h3f79840d : _GEN_146; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_148 = 11'h94 == io_cosIndex[10:0] ? 30'h3f796d7d : _GEN_147; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_149 = 11'h95 == io_cosIndex[10:0] ? 30'h3f7956c6 : _GEN_148; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_150 = 11'h96 == io_cosIndex[10:0] ? 30'h3f793fe9 : _GEN_149; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_151 = 11'h97 == io_cosIndex[10:0] ? 30'h3f7928e5 : _GEN_150; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_152 = 11'h98 == io_cosIndex[10:0] ? 30'h3f7911bb : _GEN_151; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_153 = 11'h99 == io_cosIndex[10:0] ? 30'h3f78fa6a : _GEN_152; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_154 = 11'h9a == io_cosIndex[10:0] ? 30'h3f78e2f3 : _GEN_153; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_155 = 11'h9b == io_cosIndex[10:0] ? 30'h3f78cb56 : _GEN_154; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_156 = 11'h9c == io_cosIndex[10:0] ? 30'h3f78b392 : _GEN_155; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_157 = 11'h9d == io_cosIndex[10:0] ? 30'h3f789ba8 : _GEN_156; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_158 = 11'h9e == io_cosIndex[10:0] ? 30'h3f788398 : _GEN_157; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_159 = 11'h9f == io_cosIndex[10:0] ? 30'h3f786b61 : _GEN_158; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_160 = 11'ha0 == io_cosIndex[10:0] ? 30'h3f785304 : _GEN_159; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_161 = 11'ha1 == io_cosIndex[10:0] ? 30'h3f783a80 : _GEN_160; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_162 = 11'ha2 == io_cosIndex[10:0] ? 30'h3f7821d6 : _GEN_161; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_163 = 11'ha3 == io_cosIndex[10:0] ? 30'h3f780906 : _GEN_162; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_164 = 11'ha4 == io_cosIndex[10:0] ? 30'h3f77f010 : _GEN_163; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_165 = 11'ha5 == io_cosIndex[10:0] ? 30'h3f77d6f3 : _GEN_164; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_166 = 11'ha6 == io_cosIndex[10:0] ? 30'h3f77bdb0 : _GEN_165; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_167 = 11'ha7 == io_cosIndex[10:0] ? 30'h3f77a447 : _GEN_166; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_168 = 11'ha8 == io_cosIndex[10:0] ? 30'h3f778ab8 : _GEN_167; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_169 = 11'ha9 == io_cosIndex[10:0] ? 30'h3f777103 : _GEN_168; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_170 = 11'haa == io_cosIndex[10:0] ? 30'h3f775727 : _GEN_169; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_171 = 11'hab == io_cosIndex[10:0] ? 30'h3f773d25 : _GEN_170; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_172 = 11'hac == io_cosIndex[10:0] ? 30'h3f7722fd : _GEN_171; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_173 = 11'had == io_cosIndex[10:0] ? 30'h3f7708af : _GEN_172; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_174 = 11'hae == io_cosIndex[10:0] ? 30'h3f76ee3b : _GEN_173; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_175 = 11'haf == io_cosIndex[10:0] ? 30'h3f76d3a1 : _GEN_174; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_176 = 11'hb0 == io_cosIndex[10:0] ? 30'h3f76b8e0 : _GEN_175; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_177 = 11'hb1 == io_cosIndex[10:0] ? 30'h3f769dfa : _GEN_176; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_178 = 11'hb2 == io_cosIndex[10:0] ? 30'h3f7682ed : _GEN_177; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_179 = 11'hb3 == io_cosIndex[10:0] ? 30'h3f7667bb : _GEN_178; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_180 = 11'hb4 == io_cosIndex[10:0] ? 30'h3f764c62 : _GEN_179; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_181 = 11'hb5 == io_cosIndex[10:0] ? 30'h3f7630e4 : _GEN_180; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_182 = 11'hb6 == io_cosIndex[10:0] ? 30'h3f76153f : _GEN_181; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_183 = 11'hb7 == io_cosIndex[10:0] ? 30'h3f75f975 : _GEN_182; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_184 = 11'hb8 == io_cosIndex[10:0] ? 30'h3f75dd84 : _GEN_183; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_185 = 11'hb9 == io_cosIndex[10:0] ? 30'h3f75c16e : _GEN_184; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_186 = 11'hba == io_cosIndex[10:0] ? 30'h3f75a531 : _GEN_185; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_187 = 11'hbb == io_cosIndex[10:0] ? 30'h3f7588cf : _GEN_186; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_188 = 11'hbc == io_cosIndex[10:0] ? 30'h3f756c47 : _GEN_187; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_189 = 11'hbd == io_cosIndex[10:0] ? 30'h3f754f99 : _GEN_188; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_190 = 11'hbe == io_cosIndex[10:0] ? 30'h3f7532c5 : _GEN_189; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_191 = 11'hbf == io_cosIndex[10:0] ? 30'h3f7515cc : _GEN_190; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_192 = 11'hc0 == io_cosIndex[10:0] ? 30'h3f74f8ac : _GEN_191; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_193 = 11'hc1 == io_cosIndex[10:0] ? 30'h3f74db67 : _GEN_192; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_194 = 11'hc2 == io_cosIndex[10:0] ? 30'h3f74bdfc : _GEN_193; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_195 = 11'hc3 == io_cosIndex[10:0] ? 30'h3f74a06b : _GEN_194; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_196 = 11'hc4 == io_cosIndex[10:0] ? 30'h3f7482b5 : _GEN_195; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_197 = 11'hc5 == io_cosIndex[10:0] ? 30'h3f7464d9 : _GEN_196; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_198 = 11'hc6 == io_cosIndex[10:0] ? 30'h3f7446d7 : _GEN_197; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_199 = 11'hc7 == io_cosIndex[10:0] ? 30'h3f7428af : _GEN_198; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_200 = 11'hc8 == io_cosIndex[10:0] ? 30'h3f740a62 : _GEN_199; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_201 = 11'hc9 == io_cosIndex[10:0] ? 30'h3f73ebef : _GEN_200; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_202 = 11'hca == io_cosIndex[10:0] ? 30'h3f73cd56 : _GEN_201; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_203 = 11'hcb == io_cosIndex[10:0] ? 30'h3f73ae98 : _GEN_202; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_204 = 11'hcc == io_cosIndex[10:0] ? 30'h3f738fb4 : _GEN_203; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_205 = 11'hcd == io_cosIndex[10:0] ? 30'h3f7370ab : _GEN_204; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_206 = 11'hce == io_cosIndex[10:0] ? 30'h3f73517c : _GEN_205; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_207 = 11'hcf == io_cosIndex[10:0] ? 30'h3f733227 : _GEN_206; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_208 = 11'hd0 == io_cosIndex[10:0] ? 30'h3f7312ad : _GEN_207; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_209 = 11'hd1 == io_cosIndex[10:0] ? 30'h3f72f30e : _GEN_208; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_210 = 11'hd2 == io_cosIndex[10:0] ? 30'h3f72d349 : _GEN_209; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_211 = 11'hd3 == io_cosIndex[10:0] ? 30'h3f72b35e : _GEN_210; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_212 = 11'hd4 == io_cosIndex[10:0] ? 30'h3f72934e : _GEN_211; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_213 = 11'hd5 == io_cosIndex[10:0] ? 30'h3f727319 : _GEN_212; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_214 = 11'hd6 == io_cosIndex[10:0] ? 30'h3f7252be : _GEN_213; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_215 = 11'hd7 == io_cosIndex[10:0] ? 30'h3f72323e : _GEN_214; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_216 = 11'hd8 == io_cosIndex[10:0] ? 30'h3f721199 : _GEN_215; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_217 = 11'hd9 == io_cosIndex[10:0] ? 30'h3f71f0ce : _GEN_216; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_218 = 11'hda == io_cosIndex[10:0] ? 30'h3f71cfde : _GEN_217; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_219 = 11'hdb == io_cosIndex[10:0] ? 30'h3f71aec8 : _GEN_218; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_220 = 11'hdc == io_cosIndex[10:0] ? 30'h3f718d8d : _GEN_219; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_221 = 11'hdd == io_cosIndex[10:0] ? 30'h3f716c2d : _GEN_220; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_222 = 11'hde == io_cosIndex[10:0] ? 30'h3f714aa8 : _GEN_221; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_223 = 11'hdf == io_cosIndex[10:0] ? 30'h3f7128fe : _GEN_222; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_224 = 11'he0 == io_cosIndex[10:0] ? 30'h3f71072e : _GEN_223; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_225 = 11'he1 == io_cosIndex[10:0] ? 30'h3f70e539 : _GEN_224; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_226 = 11'he2 == io_cosIndex[10:0] ? 30'h3f70c31f : _GEN_225; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_227 = 11'he3 == io_cosIndex[10:0] ? 30'h3f70a0e0 : _GEN_226; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_228 = 11'he4 == io_cosIndex[10:0] ? 30'h3f707e7b : _GEN_227; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_229 = 11'he5 == io_cosIndex[10:0] ? 30'h3f705bf2 : _GEN_228; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_230 = 11'he6 == io_cosIndex[10:0] ? 30'h3f703943 : _GEN_229; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_231 = 11'he7 == io_cosIndex[10:0] ? 30'h3f701670 : _GEN_230; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_232 = 11'he8 == io_cosIndex[10:0] ? 30'h3f6ff377 : _GEN_231; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_233 = 11'he9 == io_cosIndex[10:0] ? 30'h3f6fd059 : _GEN_232; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_234 = 11'hea == io_cosIndex[10:0] ? 30'h3f6fad17 : _GEN_233; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_235 = 11'heb == io_cosIndex[10:0] ? 30'h3f6f89af : _GEN_234; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_236 = 11'hec == io_cosIndex[10:0] ? 30'h3f6f6622 : _GEN_235; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_237 = 11'hed == io_cosIndex[10:0] ? 30'h3f6f4271 : _GEN_236; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_238 = 11'hee == io_cosIndex[10:0] ? 30'h3f6f1e9a : _GEN_237; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_239 = 11'hef == io_cosIndex[10:0] ? 30'h3f6efa9f : _GEN_238; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_240 = 11'hf0 == io_cosIndex[10:0] ? 30'h3f6ed67f : _GEN_239; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_241 = 11'hf1 == io_cosIndex[10:0] ? 30'h3f6eb23a : _GEN_240; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_242 = 11'hf2 == io_cosIndex[10:0] ? 30'h3f6e8dd0 : _GEN_241; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_243 = 11'hf3 == io_cosIndex[10:0] ? 30'h3f6e6941 : _GEN_242; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_244 = 11'hf4 == io_cosIndex[10:0] ? 30'h3f6e448e : _GEN_243; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_245 = 11'hf5 == io_cosIndex[10:0] ? 30'h3f6e1fb5 : _GEN_244; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_246 = 11'hf6 == io_cosIndex[10:0] ? 30'h3f6dfab8 : _GEN_245; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_247 = 11'hf7 == io_cosIndex[10:0] ? 30'h3f6dd597 : _GEN_246; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_248 = 11'hf8 == io_cosIndex[10:0] ? 30'h3f6db050 : _GEN_247; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_249 = 11'hf9 == io_cosIndex[10:0] ? 30'h3f6d8ae5 : _GEN_248; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_250 = 11'hfa == io_cosIndex[10:0] ? 30'h3f6d6555 : _GEN_249; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_251 = 11'hfb == io_cosIndex[10:0] ? 30'h3f6d3fa1 : _GEN_250; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_252 = 11'hfc == io_cosIndex[10:0] ? 30'h3f6d19c8 : _GEN_251; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_253 = 11'hfd == io_cosIndex[10:0] ? 30'h3f6cf3cb : _GEN_252; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_254 = 11'hfe == io_cosIndex[10:0] ? 30'h3f6ccda8 : _GEN_253; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_255 = 11'hff == io_cosIndex[10:0] ? 30'h3f6ca762 : _GEN_254; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_256 = 11'h100 == io_cosIndex[10:0] ? 30'h3f6c80f7 : _GEN_255; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_257 = 11'h101 == io_cosIndex[10:0] ? 30'h3f6c5a67 : _GEN_256; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_258 = 11'h102 == io_cosIndex[10:0] ? 30'h3f6c33b3 : _GEN_257; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_259 = 11'h103 == io_cosIndex[10:0] ? 30'h3f6c0cda : _GEN_258; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_260 = 11'h104 == io_cosIndex[10:0] ? 30'h3f6be5dd : _GEN_259; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_261 = 11'h105 == io_cosIndex[10:0] ? 30'h3f6bbebc : _GEN_260; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_262 = 11'h106 == io_cosIndex[10:0] ? 30'h3f6b9776 : _GEN_261; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_263 = 11'h107 == io_cosIndex[10:0] ? 30'h3f6b700c : _GEN_262; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_264 = 11'h108 == io_cosIndex[10:0] ? 30'h3f6b487e : _GEN_263; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_265 = 11'h109 == io_cosIndex[10:0] ? 30'h3f6b20cb : _GEN_264; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_266 = 11'h10a == io_cosIndex[10:0] ? 30'h3f6af8f4 : _GEN_265; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_267 = 11'h10b == io_cosIndex[10:0] ? 30'h3f6ad0f9 : _GEN_266; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_268 = 11'h10c == io_cosIndex[10:0] ? 30'h3f6aa8d9 : _GEN_267; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_269 = 11'h10d == io_cosIndex[10:0] ? 30'h3f6a8096 : _GEN_268; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_270 = 11'h10e == io_cosIndex[10:0] ? 30'h3f6a582e : _GEN_269; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_271 = 11'h10f == io_cosIndex[10:0] ? 30'h3f6a2fa2 : _GEN_270; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_272 = 11'h110 == io_cosIndex[10:0] ? 30'h3f6a06f2 : _GEN_271; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_273 = 11'h111 == io_cosIndex[10:0] ? 30'h3f69de1d : _GEN_272; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_274 = 11'h112 == io_cosIndex[10:0] ? 30'h3f69b525 : _GEN_273; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_275 = 11'h113 == io_cosIndex[10:0] ? 30'h3f698c09 : _GEN_274; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_276 = 11'h114 == io_cosIndex[10:0] ? 30'h3f6962c8 : _GEN_275; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_277 = 11'h115 == io_cosIndex[10:0] ? 30'h3f693964 : _GEN_276; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_278 = 11'h116 == io_cosIndex[10:0] ? 30'h3f690fdb : _GEN_277; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_279 = 11'h117 == io_cosIndex[10:0] ? 30'h3f68e62f : _GEN_278; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_280 = 11'h118 == io_cosIndex[10:0] ? 30'h3f68bc5f : _GEN_279; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_281 = 11'h119 == io_cosIndex[10:0] ? 30'h3f68926b : _GEN_280; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_282 = 11'h11a == io_cosIndex[10:0] ? 30'h3f686852 : _GEN_281; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_283 = 11'h11b == io_cosIndex[10:0] ? 30'h3f683e16 : _GEN_282; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_284 = 11'h11c == io_cosIndex[10:0] ? 30'h3f6813b7 : _GEN_283; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_285 = 11'h11d == io_cosIndex[10:0] ? 30'h3f67e933 : _GEN_284; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_286 = 11'h11e == io_cosIndex[10:0] ? 30'h3f67be8c : _GEN_285; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_287 = 11'h11f == io_cosIndex[10:0] ? 30'h3f6793c1 : _GEN_286; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_288 = 11'h120 == io_cosIndex[10:0] ? 30'h3f6768d2 : _GEN_287; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_289 = 11'h121 == io_cosIndex[10:0] ? 30'h3f673dbf : _GEN_288; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_290 = 11'h122 == io_cosIndex[10:0] ? 30'h3f671289 : _GEN_289; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_291 = 11'h123 == io_cosIndex[10:0] ? 30'h3f66e72f : _GEN_290; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_292 = 11'h124 == io_cosIndex[10:0] ? 30'h3f66bbb1 : _GEN_291; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_293 = 11'h125 == io_cosIndex[10:0] ? 30'h3f669010 : _GEN_292; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_294 = 11'h126 == io_cosIndex[10:0] ? 30'h3f66644c : _GEN_293; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_295 = 11'h127 == io_cosIndex[10:0] ? 30'h3f663863 : _GEN_294; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_296 = 11'h128 == io_cosIndex[10:0] ? 30'h3f660c58 : _GEN_295; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_297 = 11'h129 == io_cosIndex[10:0] ? 30'h3f65e028 : _GEN_296; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_298 = 11'h12a == io_cosIndex[10:0] ? 30'h3f65b3d6 : _GEN_297; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_299 = 11'h12b == io_cosIndex[10:0] ? 30'h3f65875f : _GEN_298; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_300 = 11'h12c == io_cosIndex[10:0] ? 30'h3f655ac6 : _GEN_299; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_301 = 11'h12d == io_cosIndex[10:0] ? 30'h3f652e09 : _GEN_300; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_302 = 11'h12e == io_cosIndex[10:0] ? 30'h3f650129 : _GEN_301; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_303 = 11'h12f == io_cosIndex[10:0] ? 30'h3f64d425 : _GEN_302; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_304 = 11'h130 == io_cosIndex[10:0] ? 30'h3f64a6fe : _GEN_303; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_305 = 11'h131 == io_cosIndex[10:0] ? 30'h3f6479b4 : _GEN_304; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_306 = 11'h132 == io_cosIndex[10:0] ? 30'h3f644c46 : _GEN_305; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_307 = 11'h133 == io_cosIndex[10:0] ? 30'h3f641eb5 : _GEN_306; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_308 = 11'h134 == io_cosIndex[10:0] ? 30'h3f63f102 : _GEN_307; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_309 = 11'h135 == io_cosIndex[10:0] ? 30'h3f63c32a : _GEN_308; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_310 = 11'h136 == io_cosIndex[10:0] ? 30'h3f639530 : _GEN_309; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_311 = 11'h137 == io_cosIndex[10:0] ? 30'h3f636713 : _GEN_310; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_312 = 11'h138 == io_cosIndex[10:0] ? 30'h3f6338d3 : _GEN_311; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_313 = 11'h139 == io_cosIndex[10:0] ? 30'h3f630a6f : _GEN_312; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_314 = 11'h13a == io_cosIndex[10:0] ? 30'h3f62dbe9 : _GEN_313; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_315 = 11'h13b == io_cosIndex[10:0] ? 30'h3f62ad3f : _GEN_314; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_316 = 11'h13c == io_cosIndex[10:0] ? 30'h3f627e73 : _GEN_315; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_317 = 11'h13d == io_cosIndex[10:0] ? 30'h3f624f83 : _GEN_316; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_318 = 11'h13e == io_cosIndex[10:0] ? 30'h3f622071 : _GEN_317; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_319 = 11'h13f == io_cosIndex[10:0] ? 30'h3f61f13c : _GEN_318; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_320 = 11'h140 == io_cosIndex[10:0] ? 30'h3f61c1e3 : _GEN_319; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_321 = 11'h141 == io_cosIndex[10:0] ? 30'h3f619268 : _GEN_320; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_322 = 11'h142 == io_cosIndex[10:0] ? 30'h3f6162cb : _GEN_321; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_323 = 11'h143 == io_cosIndex[10:0] ? 30'h3f61330a : _GEN_322; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_324 = 11'h144 == io_cosIndex[10:0] ? 30'h3f610327 : _GEN_323; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_325 = 11'h145 == io_cosIndex[10:0] ? 30'h3f60d321 : _GEN_324; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_326 = 11'h146 == io_cosIndex[10:0] ? 30'h3f60a2f8 : _GEN_325; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_327 = 11'h147 == io_cosIndex[10:0] ? 30'h3f6072ad : _GEN_326; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_328 = 11'h148 == io_cosIndex[10:0] ? 30'h3f60423f : _GEN_327; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_329 = 11'h149 == io_cosIndex[10:0] ? 30'h3f6011af : _GEN_328; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_330 = 11'h14a == io_cosIndex[10:0] ? 30'h3f5fe0fb : _GEN_329; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_331 = 11'h14b == io_cosIndex[10:0] ? 30'h3f5fb026 : _GEN_330; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_332 = 11'h14c == io_cosIndex[10:0] ? 30'h3f5f7f2e : _GEN_331; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_333 = 11'h14d == io_cosIndex[10:0] ? 30'h3f5f4e13 : _GEN_332; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_334 = 11'h14e == io_cosIndex[10:0] ? 30'h3f5f1cd6 : _GEN_333; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_335 = 11'h14f == io_cosIndex[10:0] ? 30'h3f5eeb76 : _GEN_334; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_336 = 11'h150 == io_cosIndex[10:0] ? 30'h3f5eb9f4 : _GEN_335; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_337 = 11'h151 == io_cosIndex[10:0] ? 30'h3f5e8850 : _GEN_336; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_338 = 11'h152 == io_cosIndex[10:0] ? 30'h3f5e568a : _GEN_337; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_339 = 11'h153 == io_cosIndex[10:0] ? 30'h3f5e24a1 : _GEN_338; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_340 = 11'h154 == io_cosIndex[10:0] ? 30'h3f5df295 : _GEN_339; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_341 = 11'h155 == io_cosIndex[10:0] ? 30'h3f5dc068 : _GEN_340; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_342 = 11'h156 == io_cosIndex[10:0] ? 30'h3f5d8e18 : _GEN_341; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_343 = 11'h157 == io_cosIndex[10:0] ? 30'h3f5d5ba6 : _GEN_342; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_344 = 11'h158 == io_cosIndex[10:0] ? 30'h3f5d2912 : _GEN_343; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_345 = 11'h159 == io_cosIndex[10:0] ? 30'h3f5cf65c : _GEN_344; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_346 = 11'h15a == io_cosIndex[10:0] ? 30'h3f5cc384 : _GEN_345; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_347 = 11'h15b == io_cosIndex[10:0] ? 30'h3f5c908a : _GEN_346; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_348 = 11'h15c == io_cosIndex[10:0] ? 30'h3f5c5d6e : _GEN_347; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_349 = 11'h15d == io_cosIndex[10:0] ? 30'h3f5c2a2f : _GEN_348; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_350 = 11'h15e == io_cosIndex[10:0] ? 30'h3f5bf6cf : _GEN_349; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_351 = 11'h15f == io_cosIndex[10:0] ? 30'h3f5bc34d : _GEN_350; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_352 = 11'h160 == io_cosIndex[10:0] ? 30'h3f5b8fa9 : _GEN_351; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_353 = 11'h161 == io_cosIndex[10:0] ? 30'h3f5b5be3 : _GEN_352; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_354 = 11'h162 == io_cosIndex[10:0] ? 30'h3f5b27fb : _GEN_353; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_355 = 11'h163 == io_cosIndex[10:0] ? 30'h3f5af3f1 : _GEN_354; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_356 = 11'h164 == io_cosIndex[10:0] ? 30'h3f5abfc6 : _GEN_355; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_357 = 11'h165 == io_cosIndex[10:0] ? 30'h3f5a8b79 : _GEN_356; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_358 = 11'h166 == io_cosIndex[10:0] ? 30'h3f5a570a : _GEN_357; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_359 = 11'h167 == io_cosIndex[10:0] ? 30'h3f5a2279 : _GEN_358; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_360 = 11'h168 == io_cosIndex[10:0] ? 30'h3f59edc7 : _GEN_359; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_361 = 11'h169 == io_cosIndex[10:0] ? 30'h3f59b8f3 : _GEN_360; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_362 = 11'h16a == io_cosIndex[10:0] ? 30'h3f5983fe : _GEN_361; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_363 = 11'h16b == io_cosIndex[10:0] ? 30'h3f594ee7 : _GEN_362; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_364 = 11'h16c == io_cosIndex[10:0] ? 30'h3f5919ae : _GEN_363; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_365 = 11'h16d == io_cosIndex[10:0] ? 30'h3f58e454 : _GEN_364; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_366 = 11'h16e == io_cosIndex[10:0] ? 30'h3f58aed9 : _GEN_365; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_367 = 11'h16f == io_cosIndex[10:0] ? 30'h3f58793c : _GEN_366; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_368 = 11'h170 == io_cosIndex[10:0] ? 30'h3f58437d : _GEN_367; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_369 = 11'h171 == io_cosIndex[10:0] ? 30'h3f580d9e : _GEN_368; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_370 = 11'h172 == io_cosIndex[10:0] ? 30'h3f57d79d : _GEN_369; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_371 = 11'h173 == io_cosIndex[10:0] ? 30'h3f57a17a : _GEN_370; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_372 = 11'h174 == io_cosIndex[10:0] ? 30'h3f576b37 : _GEN_371; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_373 = 11'h175 == io_cosIndex[10:0] ? 30'h3f5734d2 : _GEN_372; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_374 = 11'h176 == io_cosIndex[10:0] ? 30'h3f56fe4c : _GEN_373; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_375 = 11'h177 == io_cosIndex[10:0] ? 30'h3f56c7a5 : _GEN_374; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_376 = 11'h178 == io_cosIndex[10:0] ? 30'h3f5690dc : _GEN_375; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_377 = 11'h179 == io_cosIndex[10:0] ? 30'h3f5659f3 : _GEN_376; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_378 = 11'h17a == io_cosIndex[10:0] ? 30'h3f5622e8 : _GEN_377; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_379 = 11'h17b == io_cosIndex[10:0] ? 30'h3f55ebbd : _GEN_378; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_380 = 11'h17c == io_cosIndex[10:0] ? 30'h3f55b470 : _GEN_379; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_381 = 11'h17d == io_cosIndex[10:0] ? 30'h3f557d02 : _GEN_380; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_382 = 11'h17e == io_cosIndex[10:0] ? 30'h3f554574 : _GEN_381; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_383 = 11'h17f == io_cosIndex[10:0] ? 30'h3f550dc5 : _GEN_382; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_384 = 11'h180 == io_cosIndex[10:0] ? 30'h3f54d5f4 : _GEN_383; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_385 = 11'h181 == io_cosIndex[10:0] ? 30'h3f549e03 : _GEN_384; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_386 = 11'h182 == io_cosIndex[10:0] ? 30'h3f5465f1 : _GEN_385; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_387 = 11'h183 == io_cosIndex[10:0] ? 30'h3f542dbf : _GEN_386; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_388 = 11'h184 == io_cosIndex[10:0] ? 30'h3f53f56b : _GEN_387; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_389 = 11'h185 == io_cosIndex[10:0] ? 30'h3f53bcf7 : _GEN_388; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_390 = 11'h186 == io_cosIndex[10:0] ? 30'h3f538462 : _GEN_389; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_391 = 11'h187 == io_cosIndex[10:0] ? 30'h3f534bad : _GEN_390; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_392 = 11'h188 == io_cosIndex[10:0] ? 30'h3f5312d7 : _GEN_391; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_393 = 11'h189 == io_cosIndex[10:0] ? 30'h3f52d9e0 : _GEN_392; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_394 = 11'h18a == io_cosIndex[10:0] ? 30'h3f52a0c9 : _GEN_393; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_395 = 11'h18b == io_cosIndex[10:0] ? 30'h3f526792 : _GEN_394; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_396 = 11'h18c == io_cosIndex[10:0] ? 30'h3f522e3a : _GEN_395; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_397 = 11'h18d == io_cosIndex[10:0] ? 30'h3f51f4c1 : _GEN_396; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_398 = 11'h18e == io_cosIndex[10:0] ? 30'h3f51bb28 : _GEN_397; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_399 = 11'h18f == io_cosIndex[10:0] ? 30'h3f51816f : _GEN_398; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_400 = 11'h190 == io_cosIndex[10:0] ? 30'h3f514795 : _GEN_399; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_401 = 11'h191 == io_cosIndex[10:0] ? 30'h3f510d9b : _GEN_400; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_402 = 11'h192 == io_cosIndex[10:0] ? 30'h3f50d381 : _GEN_401; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_403 = 11'h193 == io_cosIndex[10:0] ? 30'h3f509947 : _GEN_402; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_404 = 11'h194 == io_cosIndex[10:0] ? 30'h3f505eec : _GEN_403; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_405 = 11'h195 == io_cosIndex[10:0] ? 30'h3f502472 : _GEN_404; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_406 = 11'h196 == io_cosIndex[10:0] ? 30'h3f4fe9d7 : _GEN_405; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_407 = 11'h197 == io_cosIndex[10:0] ? 30'h3f4faf1c : _GEN_406; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_408 = 11'h198 == io_cosIndex[10:0] ? 30'h3f4f7441 : _GEN_407; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_409 = 11'h199 == io_cosIndex[10:0] ? 30'h3f4f3946 : _GEN_408; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_410 = 11'h19a == io_cosIndex[10:0] ? 30'h3f4efe2b : _GEN_409; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_411 = 11'h19b == io_cosIndex[10:0] ? 30'h3f4ec2f1 : _GEN_410; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_412 = 11'h19c == io_cosIndex[10:0] ? 30'h3f4e8796 : _GEN_411; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_413 = 11'h19d == io_cosIndex[10:0] ? 30'h3f4e4c1b : _GEN_412; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_414 = 11'h19e == io_cosIndex[10:0] ? 30'h3f4e1081 : _GEN_413; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_415 = 11'h19f == io_cosIndex[10:0] ? 30'h3f4dd4c7 : _GEN_414; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_416 = 11'h1a0 == io_cosIndex[10:0] ? 30'h3f4d98ed : _GEN_415; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_417 = 11'h1a1 == io_cosIndex[10:0] ? 30'h3f4d5cf3 : _GEN_416; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_418 = 11'h1a2 == io_cosIndex[10:0] ? 30'h3f4d20da : _GEN_417; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_419 = 11'h1a3 == io_cosIndex[10:0] ? 30'h3f4ce4a1 : _GEN_418; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_420 = 11'h1a4 == io_cosIndex[10:0] ? 30'h3f4ca848 : _GEN_419; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_421 = 11'h1a5 == io_cosIndex[10:0] ? 30'h3f4c6bd0 : _GEN_420; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_422 = 11'h1a6 == io_cosIndex[10:0] ? 30'h3f4c2f38 : _GEN_421; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_423 = 11'h1a7 == io_cosIndex[10:0] ? 30'h3f4bf281 : _GEN_422; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_424 = 11'h1a8 == io_cosIndex[10:0] ? 30'h3f4bb5aa : _GEN_423; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_425 = 11'h1a9 == io_cosIndex[10:0] ? 30'h3f4b78b4 : _GEN_424; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_426 = 11'h1aa == io_cosIndex[10:0] ? 30'h3f4b3b9e : _GEN_425; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_427 = 11'h1ab == io_cosIndex[10:0] ? 30'h3f4afe69 : _GEN_426; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_428 = 11'h1ac == io_cosIndex[10:0] ? 30'h3f4ac115 : _GEN_427; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_429 = 11'h1ad == io_cosIndex[10:0] ? 30'h3f4a83a2 : _GEN_428; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_430 = 11'h1ae == io_cosIndex[10:0] ? 30'h3f4a460f : _GEN_429; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_431 = 11'h1af == io_cosIndex[10:0] ? 30'h3f4a085d : _GEN_430; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_432 = 11'h1b0 == io_cosIndex[10:0] ? 30'h3f49ca8c : _GEN_431; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_433 = 11'h1b1 == io_cosIndex[10:0] ? 30'h3f498c9c : _GEN_432; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_434 = 11'h1b2 == io_cosIndex[10:0] ? 30'h3f494e8c : _GEN_433; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_435 = 11'h1b3 == io_cosIndex[10:0] ? 30'h3f49105e : _GEN_434; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_436 = 11'h1b4 == io_cosIndex[10:0] ? 30'h3f48d210 : _GEN_435; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_437 = 11'h1b5 == io_cosIndex[10:0] ? 30'h3f4893a4 : _GEN_436; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_438 = 11'h1b6 == io_cosIndex[10:0] ? 30'h3f485518 : _GEN_437; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_439 = 11'h1b7 == io_cosIndex[10:0] ? 30'h3f48166e : _GEN_438; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_440 = 11'h1b8 == io_cosIndex[10:0] ? 30'h3f47d7a5 : _GEN_439; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_441 = 11'h1b9 == io_cosIndex[10:0] ? 30'h3f4798bd : _GEN_440; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_442 = 11'h1ba == io_cosIndex[10:0] ? 30'h3f4759b6 : _GEN_441; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_443 = 11'h1bb == io_cosIndex[10:0] ? 30'h3f471a91 : _GEN_442; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_444 = 11'h1bc == io_cosIndex[10:0] ? 30'h3f46db4c : _GEN_443; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_445 = 11'h1bd == io_cosIndex[10:0] ? 30'h3f469bea : _GEN_444; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_446 = 11'h1be == io_cosIndex[10:0] ? 30'h3f465c68 : _GEN_445; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_447 = 11'h1bf == io_cosIndex[10:0] ? 30'h3f461cc8 : _GEN_446; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_448 = 11'h1c0 == io_cosIndex[10:0] ? 30'h3f45dd09 : _GEN_447; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_449 = 11'h1c1 == io_cosIndex[10:0] ? 30'h3f459d2c : _GEN_448; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_450 = 11'h1c2 == io_cosIndex[10:0] ? 30'h3f455d30 : _GEN_449; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_451 = 11'h1c3 == io_cosIndex[10:0] ? 30'h3f451d16 : _GEN_450; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_452 = 11'h1c4 == io_cosIndex[10:0] ? 30'h3f44dcdd : _GEN_451; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_453 = 11'h1c5 == io_cosIndex[10:0] ? 30'h3f449c86 : _GEN_452; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_454 = 11'h1c6 == io_cosIndex[10:0] ? 30'h3f445c11 : _GEN_453; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_455 = 11'h1c7 == io_cosIndex[10:0] ? 30'h3f441b7d : _GEN_454; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_456 = 11'h1c8 == io_cosIndex[10:0] ? 30'h3f43dacb : _GEN_455; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_457 = 11'h1c9 == io_cosIndex[10:0] ? 30'h3f4399fb : _GEN_456; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_458 = 11'h1ca == io_cosIndex[10:0] ? 30'h3f43590d : _GEN_457; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_459 = 11'h1cb == io_cosIndex[10:0] ? 30'h3f431800 : _GEN_458; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_460 = 11'h1cc == io_cosIndex[10:0] ? 30'h3f42d6d6 : _GEN_459; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_461 = 11'h1cd == io_cosIndex[10:0] ? 30'h3f42958d : _GEN_460; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_462 = 11'h1ce == io_cosIndex[10:0] ? 30'h3f425427 : _GEN_461; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_463 = 11'h1cf == io_cosIndex[10:0] ? 30'h3f4212a2 : _GEN_462; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_464 = 11'h1d0 == io_cosIndex[10:0] ? 30'h3f41d0ff : _GEN_463; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_465 = 11'h1d1 == io_cosIndex[10:0] ? 30'h3f418f3f : _GEN_464; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_466 = 11'h1d2 == io_cosIndex[10:0] ? 30'h3f414d61 : _GEN_465; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_467 = 11'h1d3 == io_cosIndex[10:0] ? 30'h3f410b65 : _GEN_466; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_468 = 11'h1d4 == io_cosIndex[10:0] ? 30'h3f40c94b : _GEN_467; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_469 = 11'h1d5 == io_cosIndex[10:0] ? 30'h3f408713 : _GEN_468; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_470 = 11'h1d6 == io_cosIndex[10:0] ? 30'h3f4044be : _GEN_469; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_471 = 11'h1d7 == io_cosIndex[10:0] ? 30'h3f40024b : _GEN_470; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_472 = 11'h1d8 == io_cosIndex[10:0] ? 30'h3f3fbfba : _GEN_471; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_473 = 11'h1d9 == io_cosIndex[10:0] ? 30'h3f3f7d0c : _GEN_472; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_474 = 11'h1da == io_cosIndex[10:0] ? 30'h3f3f3a40 : _GEN_473; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_475 = 11'h1db == io_cosIndex[10:0] ? 30'h3f3ef757 : _GEN_474; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_476 = 11'h1dc == io_cosIndex[10:0] ? 30'h3f3eb450 : _GEN_475; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_477 = 11'h1dd == io_cosIndex[10:0] ? 30'h3f3e712c : _GEN_476; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_478 = 11'h1de == io_cosIndex[10:0] ? 30'h3f3e2dea : _GEN_477; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_479 = 11'h1df == io_cosIndex[10:0] ? 30'h3f3dea8b : _GEN_478; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_480 = 11'h1e0 == io_cosIndex[10:0] ? 30'h3f3da70f : _GEN_479; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_481 = 11'h1e1 == io_cosIndex[10:0] ? 30'h3f3d6376 : _GEN_480; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_482 = 11'h1e2 == io_cosIndex[10:0] ? 30'h3f3d1fbf : _GEN_481; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_483 = 11'h1e3 == io_cosIndex[10:0] ? 30'h3f3cdbeb : _GEN_482; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_484 = 11'h1e4 == io_cosIndex[10:0] ? 30'h3f3c97fa : _GEN_483; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_485 = 11'h1e5 == io_cosIndex[10:0] ? 30'h3f3c53ec : _GEN_484; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_486 = 11'h1e6 == io_cosIndex[10:0] ? 30'h3f3c0fc1 : _GEN_485; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_487 = 11'h1e7 == io_cosIndex[10:0] ? 30'h3f3bcb79 : _GEN_486; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_488 = 11'h1e8 == io_cosIndex[10:0] ? 30'h3f3b8713 : _GEN_487; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_489 = 11'h1e9 == io_cosIndex[10:0] ? 30'h3f3b4291 : _GEN_488; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_490 = 11'h1ea == io_cosIndex[10:0] ? 30'h3f3afdf2 : _GEN_489; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_491 = 11'h1eb == io_cosIndex[10:0] ? 30'h3f3ab937 : _GEN_490; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_492 = 11'h1ec == io_cosIndex[10:0] ? 30'h3f3a745e : _GEN_491; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_493 = 11'h1ed == io_cosIndex[10:0] ? 30'h3f3a2f68 : _GEN_492; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_494 = 11'h1ee == io_cosIndex[10:0] ? 30'h3f39ea56 : _GEN_493; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_495 = 11'h1ef == io_cosIndex[10:0] ? 30'h3f39a528 : _GEN_494; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_496 = 11'h1f0 == io_cosIndex[10:0] ? 30'h3f395fdc : _GEN_495; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_497 = 11'h1f1 == io_cosIndex[10:0] ? 30'h3f391a74 : _GEN_496; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_498 = 11'h1f2 == io_cosIndex[10:0] ? 30'h3f38d4ef : _GEN_497; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_499 = 11'h1f3 == io_cosIndex[10:0] ? 30'h3f388f4e : _GEN_498; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_500 = 11'h1f4 == io_cosIndex[10:0] ? 30'h3f384991 : _GEN_499; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_501 = 11'h1f5 == io_cosIndex[10:0] ? 30'h3f3803b7 : _GEN_500; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_502 = 11'h1f6 == io_cosIndex[10:0] ? 30'h3f37bdc0 : _GEN_501; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_503 = 11'h1f7 == io_cosIndex[10:0] ? 30'h3f3777ad : _GEN_502; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_504 = 11'h1f8 == io_cosIndex[10:0] ? 30'h3f37317e : _GEN_503; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_505 = 11'h1f9 == io_cosIndex[10:0] ? 30'h3f36eb33 : _GEN_504; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_506 = 11'h1fa == io_cosIndex[10:0] ? 30'h3f36a4cb : _GEN_505; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_507 = 11'h1fb == io_cosIndex[10:0] ? 30'h3f365e48 : _GEN_506; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_508 = 11'h1fc == io_cosIndex[10:0] ? 30'h3f3617a8 : _GEN_507; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_509 = 11'h1fd == io_cosIndex[10:0] ? 30'h3f35d0ec : _GEN_508; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_510 = 11'h1fe == io_cosIndex[10:0] ? 30'h3f358a14 : _GEN_509; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_511 = 11'h1ff == io_cosIndex[10:0] ? 30'h3f354320 : _GEN_510; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_512 = 11'h200 == io_cosIndex[10:0] ? 30'h3f34fc10 : _GEN_511; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_513 = 11'h201 == io_cosIndex[10:0] ? 30'h3f34b4e4 : _GEN_512; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_514 = 11'h202 == io_cosIndex[10:0] ? 30'h3f346d9c : _GEN_513; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_515 = 11'h203 == io_cosIndex[10:0] ? 30'h3f342638 : _GEN_514; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_516 = 11'h204 == io_cosIndex[10:0] ? 30'h3f33deb9 : _GEN_515; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_517 = 11'h205 == io_cosIndex[10:0] ? 30'h3f33971e : _GEN_516; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_518 = 11'h206 == io_cosIndex[10:0] ? 30'h3f334f67 : _GEN_517; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_519 = 11'h207 == io_cosIndex[10:0] ? 30'h3f330794 : _GEN_518; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_520 = 11'h208 == io_cosIndex[10:0] ? 30'h3f32bfa6 : _GEN_519; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_521 = 11'h209 == io_cosIndex[10:0] ? 30'h3f32779c : _GEN_520; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_522 = 11'h20a == io_cosIndex[10:0] ? 30'h3f322f77 : _GEN_521; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_523 = 11'h20b == io_cosIndex[10:0] ? 30'h3f31e736 : _GEN_522; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_524 = 11'h20c == io_cosIndex[10:0] ? 30'h3f319eda : _GEN_523; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_525 = 11'h20d == io_cosIndex[10:0] ? 30'h3f315662 : _GEN_524; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_526 = 11'h20e == io_cosIndex[10:0] ? 30'h3f310dcf : _GEN_525; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_527 = 11'h20f == io_cosIndex[10:0] ? 30'h3f30c521 : _GEN_526; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_528 = 11'h210 == io_cosIndex[10:0] ? 30'h3f307c57 : _GEN_527; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_529 = 11'h211 == io_cosIndex[10:0] ? 30'h3f303372 : _GEN_528; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_530 = 11'h212 == io_cosIndex[10:0] ? 30'h3f2fea72 : _GEN_529; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_531 = 11'h213 == io_cosIndex[10:0] ? 30'h3f2fa157 : _GEN_530; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_532 = 11'h214 == io_cosIndex[10:0] ? 30'h3f2f5821 : _GEN_531; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_533 = 11'h215 == io_cosIndex[10:0] ? 30'h3f2f0ed0 : _GEN_532; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_534 = 11'h216 == io_cosIndex[10:0] ? 30'h3f2ec563 : _GEN_533; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_535 = 11'h217 == io_cosIndex[10:0] ? 30'h3f2e7bdc : _GEN_534; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_536 = 11'h218 == io_cosIndex[10:0] ? 30'h3f2e323a : _GEN_535; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_537 = 11'h219 == io_cosIndex[10:0] ? 30'h3f2de87d : _GEN_536; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_538 = 11'h21a == io_cosIndex[10:0] ? 30'h3f2d9ea5 : _GEN_537; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_539 = 11'h21b == io_cosIndex[10:0] ? 30'h3f2d54b2 : _GEN_538; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_540 = 11'h21c == io_cosIndex[10:0] ? 30'h3f2d0aa5 : _GEN_539; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_541 = 11'h21d == io_cosIndex[10:0] ? 30'h3f2cc07c : _GEN_540; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_542 = 11'h21e == io_cosIndex[10:0] ? 30'h3f2c763a : _GEN_541; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_543 = 11'h21f == io_cosIndex[10:0] ? 30'h3f2c2bdc : _GEN_542; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_544 = 11'h220 == io_cosIndex[10:0] ? 30'h3f2be164 : _GEN_543; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_545 = 11'h221 == io_cosIndex[10:0] ? 30'h3f2b96d2 : _GEN_544; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_546 = 11'h222 == io_cosIndex[10:0] ? 30'h3f2b4c25 : _GEN_545; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_547 = 11'h223 == io_cosIndex[10:0] ? 30'h3f2b015d : _GEN_546; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_548 = 11'h224 == io_cosIndex[10:0] ? 30'h3f2ab67c : _GEN_547; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_549 = 11'h225 == io_cosIndex[10:0] ? 30'h3f2a6b7f : _GEN_548; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_550 = 11'h226 == io_cosIndex[10:0] ? 30'h3f2a2069 : _GEN_549; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_551 = 11'h227 == io_cosIndex[10:0] ? 30'h3f29d538 : _GEN_550; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_552 = 11'h228 == io_cosIndex[10:0] ? 30'h3f2989ed : _GEN_551; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_553 = 11'h229 == io_cosIndex[10:0] ? 30'h3f293e88 : _GEN_552; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_554 = 11'h22a == io_cosIndex[10:0] ? 30'h3f28f309 : _GEN_553; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_555 = 11'h22b == io_cosIndex[10:0] ? 30'h3f28a770 : _GEN_554; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_556 = 11'h22c == io_cosIndex[10:0] ? 30'h3f285bbd : _GEN_555; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_557 = 11'h22d == io_cosIndex[10:0] ? 30'h3f280ff0 : _GEN_556; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_558 = 11'h22e == io_cosIndex[10:0] ? 30'h3f27c409 : _GEN_557; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_559 = 11'h22f == io_cosIndex[10:0] ? 30'h3f277808 : _GEN_558; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_560 = 11'h230 == io_cosIndex[10:0] ? 30'h3f272bed : _GEN_559; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_561 = 11'h231 == io_cosIndex[10:0] ? 30'h3f26dfb8 : _GEN_560; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_562 = 11'h232 == io_cosIndex[10:0] ? 30'h3f26936a : _GEN_561; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_563 = 11'h233 == io_cosIndex[10:0] ? 30'h3f264702 : _GEN_562; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_564 = 11'h234 == io_cosIndex[10:0] ? 30'h3f25fa80 : _GEN_563; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_565 = 11'h235 == io_cosIndex[10:0] ? 30'h3f25ade4 : _GEN_564; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_566 = 11'h236 == io_cosIndex[10:0] ? 30'h3f256130 : _GEN_565; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_567 = 11'h237 == io_cosIndex[10:0] ? 30'h3f251461 : _GEN_566; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_568 = 11'h238 == io_cosIndex[10:0] ? 30'h3f24c779 : _GEN_567; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_569 = 11'h239 == io_cosIndex[10:0] ? 30'h3f247a78 : _GEN_568; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_570 = 11'h23a == io_cosIndex[10:0] ? 30'h3f242d5d : _GEN_569; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_571 = 11'h23b == io_cosIndex[10:0] ? 30'h3f23e029 : _GEN_570; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_572 = 11'h23c == io_cosIndex[10:0] ? 30'h3f2392dc : _GEN_571; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_573 = 11'h23d == io_cosIndex[10:0] ? 30'h3f234575 : _GEN_572; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_574 = 11'h23e == io_cosIndex[10:0] ? 30'h3f22f7f5 : _GEN_573; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_575 = 11'h23f == io_cosIndex[10:0] ? 30'h3f22aa5d : _GEN_574; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_576 = 11'h240 == io_cosIndex[10:0] ? 30'h3f225cab : _GEN_575; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_577 = 11'h241 == io_cosIndex[10:0] ? 30'h3f220ee0 : _GEN_576; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_578 = 11'h242 == io_cosIndex[10:0] ? 30'h3f21c0fc : _GEN_577; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_579 = 11'h243 == io_cosIndex[10:0] ? 30'h3f2172ff : _GEN_578; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_580 = 11'h244 == io_cosIndex[10:0] ? 30'h3f2124e9 : _GEN_579; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_581 = 11'h245 == io_cosIndex[10:0] ? 30'h3f20d6ba : _GEN_580; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_582 = 11'h246 == io_cosIndex[10:0] ? 30'h3f208872 : _GEN_581; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_583 = 11'h247 == io_cosIndex[10:0] ? 30'h3f203a12 : _GEN_582; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_584 = 11'h248 == io_cosIndex[10:0] ? 30'h3f1feb99 : _GEN_583; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_585 = 11'h249 == io_cosIndex[10:0] ? 30'h3f1f9d07 : _GEN_584; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_586 = 11'h24a == io_cosIndex[10:0] ? 30'h3f1f4e5d : _GEN_585; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_587 = 11'h24b == io_cosIndex[10:0] ? 30'h3f1eff9a : _GEN_586; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_588 = 11'h24c == io_cosIndex[10:0] ? 30'h3f1eb0be : _GEN_587; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_589 = 11'h24d == io_cosIndex[10:0] ? 30'h3f1e61ca : _GEN_588; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_590 = 11'h24e == io_cosIndex[10:0] ? 30'h3f1e12be : _GEN_589; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_591 = 11'h24f == io_cosIndex[10:0] ? 30'h3f1dc399 : _GEN_590; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_592 = 11'h250 == io_cosIndex[10:0] ? 30'h3f1d745c : _GEN_591; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_593 = 11'h251 == io_cosIndex[10:0] ? 30'h3f1d2507 : _GEN_592; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_594 = 11'h252 == io_cosIndex[10:0] ? 30'h3f1cd599 : _GEN_593; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_595 = 11'h253 == io_cosIndex[10:0] ? 30'h3f1c8613 : _GEN_594; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_596 = 11'h254 == io_cosIndex[10:0] ? 30'h3f1c3675 : _GEN_595; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_597 = 11'h255 == io_cosIndex[10:0] ? 30'h3f1be6bf : _GEN_596; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_598 = 11'h256 == io_cosIndex[10:0] ? 30'h3f1b96f1 : _GEN_597; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_599 = 11'h257 == io_cosIndex[10:0] ? 30'h3f1b470a : _GEN_598; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_600 = 11'h258 == io_cosIndex[10:0] ? 30'h3f1af70c : _GEN_599; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_601 = 11'h259 == io_cosIndex[10:0] ? 30'h3f1aa6f6 : _GEN_600; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_602 = 11'h25a == io_cosIndex[10:0] ? 30'h3f1a56c8 : _GEN_601; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_603 = 11'h25b == io_cosIndex[10:0] ? 30'h3f1a0683 : _GEN_602; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_604 = 11'h25c == io_cosIndex[10:0] ? 30'h3f19b625 : _GEN_603; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_605 = 11'h25d == io_cosIndex[10:0] ? 30'h3f1965b0 : _GEN_604; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_606 = 11'h25e == io_cosIndex[10:0] ? 30'h3f191523 : _GEN_605; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_607 = 11'h25f == io_cosIndex[10:0] ? 30'h3f18c47f : _GEN_606; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_608 = 11'h260 == io_cosIndex[10:0] ? 30'h3f1873c2 : _GEN_607; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_609 = 11'h261 == io_cosIndex[10:0] ? 30'h3f1822ef : _GEN_608; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_610 = 11'h262 == io_cosIndex[10:0] ? 30'h3f17d204 : _GEN_609; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_611 = 11'h263 == io_cosIndex[10:0] ? 30'h3f178101 : _GEN_610; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_612 = 11'h264 == io_cosIndex[10:0] ? 30'h3f172fe8 : _GEN_611; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_613 = 11'h265 == io_cosIndex[10:0] ? 30'h3f16deb6 : _GEN_612; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_614 = 11'h266 == io_cosIndex[10:0] ? 30'h3f168d6e : _GEN_613; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_615 = 11'h267 == io_cosIndex[10:0] ? 30'h3f163c0e : _GEN_614; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_616 = 11'h268 == io_cosIndex[10:0] ? 30'h3f15ea97 : _GEN_615; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_617 = 11'h269 == io_cosIndex[10:0] ? 30'h3f159909 : _GEN_616; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_618 = 11'h26a == io_cosIndex[10:0] ? 30'h3f154764 : _GEN_617; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_619 = 11'h26b == io_cosIndex[10:0] ? 30'h3f14f5a8 : _GEN_618; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_620 = 11'h26c == io_cosIndex[10:0] ? 30'h3f14a3d5 : _GEN_619; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_621 = 11'h26d == io_cosIndex[10:0] ? 30'h3f1451eb : _GEN_620; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_622 = 11'h26e == io_cosIndex[10:0] ? 30'h3f13ffea : _GEN_621; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_623 = 11'h26f == io_cosIndex[10:0] ? 30'h3f13add2 : _GEN_622; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_624 = 11'h270 == io_cosIndex[10:0] ? 30'h3f135ba4 : _GEN_623; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_625 = 11'h271 == io_cosIndex[10:0] ? 30'h3f13095f : _GEN_624; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_626 = 11'h272 == io_cosIndex[10:0] ? 30'h3f12b703 : _GEN_625; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_627 = 11'h273 == io_cosIndex[10:0] ? 30'h3f126490 : _GEN_626; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_628 = 11'h274 == io_cosIndex[10:0] ? 30'h3f121207 : _GEN_627; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_629 = 11'h275 == io_cosIndex[10:0] ? 30'h3f11bf67 : _GEN_628; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_630 = 11'h276 == io_cosIndex[10:0] ? 30'h3f116cb1 : _GEN_629; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_631 = 11'h277 == io_cosIndex[10:0] ? 30'h3f1119e4 : _GEN_630; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_632 = 11'h278 == io_cosIndex[10:0] ? 30'h3f10c701 : _GEN_631; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_633 = 11'h279 == io_cosIndex[10:0] ? 30'h3f107408 : _GEN_632; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_634 = 11'h27a == io_cosIndex[10:0] ? 30'h3f1020f8 : _GEN_633; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_635 = 11'h27b == io_cosIndex[10:0] ? 30'h3f0fcdd2 : _GEN_634; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_636 = 11'h27c == io_cosIndex[10:0] ? 30'h3f0f7a96 : _GEN_635; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_637 = 11'h27d == io_cosIndex[10:0] ? 30'h3f0f2744 : _GEN_636; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_638 = 11'h27e == io_cosIndex[10:0] ? 30'h3f0ed3dc : _GEN_637; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_639 = 11'h27f == io_cosIndex[10:0] ? 30'h3f0e805d : _GEN_638; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_640 = 11'h280 == io_cosIndex[10:0] ? 30'h3f0e2cc9 : _GEN_639; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_641 = 11'h281 == io_cosIndex[10:0] ? 30'h3f0dd91f : _GEN_640; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_642 = 11'h282 == io_cosIndex[10:0] ? 30'h3f0d855f : _GEN_641; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_643 = 11'h283 == io_cosIndex[10:0] ? 30'h3f0d3189 : _GEN_642; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_644 = 11'h284 == io_cosIndex[10:0] ? 30'h3f0cdd9d : _GEN_643; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_645 = 11'h285 == io_cosIndex[10:0] ? 30'h3f0c899c : _GEN_644; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_646 = 11'h286 == io_cosIndex[10:0] ? 30'h3f0c3584 : _GEN_645; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_647 = 11'h287 == io_cosIndex[10:0] ? 30'h3f0be158 : _GEN_646; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_648 = 11'h288 == io_cosIndex[10:0] ? 30'h3f0b8d15 : _GEN_647; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_649 = 11'h289 == io_cosIndex[10:0] ? 30'h3f0b38bd : _GEN_648; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_650 = 11'h28a == io_cosIndex[10:0] ? 30'h3f0ae450 : _GEN_649; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_651 = 11'h28b == io_cosIndex[10:0] ? 30'h3f0a8fcd : _GEN_650; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_652 = 11'h28c == io_cosIndex[10:0] ? 30'h3f0a3b35 : _GEN_651; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_653 = 11'h28d == io_cosIndex[10:0] ? 30'h3f09e687 : _GEN_652; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_654 = 11'h28e == io_cosIndex[10:0] ? 30'h3f0991c4 : _GEN_653; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_655 = 11'h28f == io_cosIndex[10:0] ? 30'h3f093cec : _GEN_654; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_656 = 11'h290 == io_cosIndex[10:0] ? 30'h3f08e7ff : _GEN_655; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_657 = 11'h291 == io_cosIndex[10:0] ? 30'h3f0892fd : _GEN_656; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_658 = 11'h292 == io_cosIndex[10:0] ? 30'h3f083de5 : _GEN_657; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_659 = 11'h293 == io_cosIndex[10:0] ? 30'h3f07e8b9 : _GEN_658; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_660 = 11'h294 == io_cosIndex[10:0] ? 30'h3f079378 : _GEN_659; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_661 = 11'h295 == io_cosIndex[10:0] ? 30'h3f073e21 : _GEN_660; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_662 = 11'h296 == io_cosIndex[10:0] ? 30'h3f06e8b6 : _GEN_661; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_663 = 11'h297 == io_cosIndex[10:0] ? 30'h3f069336 : _GEN_662; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_664 = 11'h298 == io_cosIndex[10:0] ? 30'h3f063da1 : _GEN_663; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_665 = 11'h299 == io_cosIndex[10:0] ? 30'h3f05e7f8 : _GEN_664; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_666 = 11'h29a == io_cosIndex[10:0] ? 30'h3f05923a : _GEN_665; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_667 = 11'h29b == io_cosIndex[10:0] ? 30'h3f053c67 : _GEN_666; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_668 = 11'h29c == io_cosIndex[10:0] ? 30'h3f04e680 : _GEN_667; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_669 = 11'h29d == io_cosIndex[10:0] ? 30'h3f049084 : _GEN_668; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_670 = 11'h29e == io_cosIndex[10:0] ? 30'h3f043a74 : _GEN_669; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_671 = 11'h29f == io_cosIndex[10:0] ? 30'h3f03e44f : _GEN_670; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_672 = 11'h2a0 == io_cosIndex[10:0] ? 30'h3f038e16 : _GEN_671; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_673 = 11'h2a1 == io_cosIndex[10:0] ? 30'h3f0337c9 : _GEN_672; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_674 = 11'h2a2 == io_cosIndex[10:0] ? 30'h3f02e167 : _GEN_673; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_675 = 11'h2a3 == io_cosIndex[10:0] ? 30'h3f028af1 : _GEN_674; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_676 = 11'h2a4 == io_cosIndex[10:0] ? 30'h3f023468 : _GEN_675; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_677 = 11'h2a5 == io_cosIndex[10:0] ? 30'h3f01ddca : _GEN_676; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_678 = 11'h2a6 == io_cosIndex[10:0] ? 30'h3f018718 : _GEN_677; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_679 = 11'h2a7 == io_cosIndex[10:0] ? 30'h3f013052 : _GEN_678; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_680 = 11'h2a8 == io_cosIndex[10:0] ? 30'h3f00d978 : _GEN_679; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_681 = 11'h2a9 == io_cosIndex[10:0] ? 30'h3f00828a : _GEN_680; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_682 = 11'h2aa == io_cosIndex[10:0] ? 30'h3f002b88 : _GEN_681; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_683 = 11'h2ab == io_cosIndex[10:0] ? 30'h3effa8e6 : _GEN_682; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_684 = 11'h2ac == io_cosIndex[10:0] ? 30'h3efefa93 : _GEN_683; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_685 = 11'h2ad == io_cosIndex[10:0] ? 30'h3efe4c1a : _GEN_684; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_686 = 11'h2ae == io_cosIndex[10:0] ? 30'h3efd9d79 : _GEN_685; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_687 = 11'h2af == io_cosIndex[10:0] ? 30'h3efceeb1 : _GEN_686; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_688 = 11'h2b0 == io_cosIndex[10:0] ? 30'h3efc3fc2 : _GEN_687; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_689 = 11'h2b1 == io_cosIndex[10:0] ? 30'h3efb90ac : _GEN_688; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_690 = 11'h2b2 == io_cosIndex[10:0] ? 30'h3efae16f : _GEN_689; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_691 = 11'h2b3 == io_cosIndex[10:0] ? 30'h3efa320c : _GEN_690; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_692 = 11'h2b4 == io_cosIndex[10:0] ? 30'h3ef98282 : _GEN_691; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_693 = 11'h2b5 == io_cosIndex[10:0] ? 30'h3ef8d2d1 : _GEN_692; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_694 = 11'h2b6 == io_cosIndex[10:0] ? 30'h3ef822fa : _GEN_693; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_695 = 11'h2b7 == io_cosIndex[10:0] ? 30'h3ef772fd : _GEN_694; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_696 = 11'h2b8 == io_cosIndex[10:0] ? 30'h3ef6c2da : _GEN_695; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_697 = 11'h2b9 == io_cosIndex[10:0] ? 30'h3ef61290 : _GEN_696; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_698 = 11'h2ba == io_cosIndex[10:0] ? 30'h3ef56221 : _GEN_697; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_699 = 11'h2bb == io_cosIndex[10:0] ? 30'h3ef4b18c : _GEN_698; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_700 = 11'h2bc == io_cosIndex[10:0] ? 30'h3ef400d1 : _GEN_699; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_701 = 11'h2bd == io_cosIndex[10:0] ? 30'h3ef34ff0 : _GEN_700; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_702 = 11'h2be == io_cosIndex[10:0] ? 30'h3ef29eea : _GEN_701; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_703 = 11'h2bf == io_cosIndex[10:0] ? 30'h3ef1edbe : _GEN_702; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_704 = 11'h2c0 == io_cosIndex[10:0] ? 30'h3ef13c6d : _GEN_703; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_705 = 11'h2c1 == io_cosIndex[10:0] ? 30'h3ef08af7 : _GEN_704; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_706 = 11'h2c2 == io_cosIndex[10:0] ? 30'h3eefd95c : _GEN_705; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_707 = 11'h2c3 == io_cosIndex[10:0] ? 30'h3eef279b : _GEN_706; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_708 = 11'h2c4 == io_cosIndex[10:0] ? 30'h3eee75b6 : _GEN_707; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_709 = 11'h2c5 == io_cosIndex[10:0] ? 30'h3eedc3ac : _GEN_708; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_710 = 11'h2c6 == io_cosIndex[10:0] ? 30'h3eed117d : _GEN_709; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_711 = 11'h2c7 == io_cosIndex[10:0] ? 30'h3eec5f2a : _GEN_710; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_712 = 11'h2c8 == io_cosIndex[10:0] ? 30'h3eebacb2 : _GEN_711; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_713 = 11'h2c9 == io_cosIndex[10:0] ? 30'h3eeafa16 : _GEN_712; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_714 = 11'h2ca == io_cosIndex[10:0] ? 30'h3eea4756 : _GEN_713; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_715 = 11'h2cb == io_cosIndex[10:0] ? 30'h3ee99471 : _GEN_714; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_716 = 11'h2cc == io_cosIndex[10:0] ? 30'h3ee8e169 : _GEN_715; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_717 = 11'h2cd == io_cosIndex[10:0] ? 30'h3ee82e3c : _GEN_716; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_718 = 11'h2ce == io_cosIndex[10:0] ? 30'h3ee77aec : _GEN_717; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_719 = 11'h2cf == io_cosIndex[10:0] ? 30'h3ee6c778 : _GEN_718; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_720 = 11'h2d0 == io_cosIndex[10:0] ? 30'h3ee613e1 : _GEN_719; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_721 = 11'h2d1 == io_cosIndex[10:0] ? 30'h3ee56025 : _GEN_720; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_722 = 11'h2d2 == io_cosIndex[10:0] ? 30'h3ee4ac47 : _GEN_721; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_723 = 11'h2d3 == io_cosIndex[10:0] ? 30'h3ee3f845 : _GEN_722; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_724 = 11'h2d4 == io_cosIndex[10:0] ? 30'h3ee34420 : _GEN_723; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_725 = 11'h2d5 == io_cosIndex[10:0] ? 30'h3ee28fd8 : _GEN_724; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_726 = 11'h2d6 == io_cosIndex[10:0] ? 30'h3ee1db6d : _GEN_725; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_727 = 11'h2d7 == io_cosIndex[10:0] ? 30'h3ee126df : _GEN_726; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_728 = 11'h2d8 == io_cosIndex[10:0] ? 30'h3ee0722f : _GEN_727; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_729 = 11'h2d9 == io_cosIndex[10:0] ? 30'h3edfbd5c : _GEN_728; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_730 = 11'h2da == io_cosIndex[10:0] ? 30'h3edf0866 : _GEN_729; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_731 = 11'h2db == io_cosIndex[10:0] ? 30'h3ede534e : _GEN_730; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_732 = 11'h2dc == io_cosIndex[10:0] ? 30'h3edd9e13 : _GEN_731; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_733 = 11'h2dd == io_cosIndex[10:0] ? 30'h3edce8b7 : _GEN_732; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_734 = 11'h2de == io_cosIndex[10:0] ? 30'h3edc3338 : _GEN_733; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_735 = 11'h2df == io_cosIndex[10:0] ? 30'h3edb7d97 : _GEN_734; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_736 = 11'h2e0 == io_cosIndex[10:0] ? 30'h3edac7d5 : _GEN_735; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_737 = 11'h2e1 == io_cosIndex[10:0] ? 30'h3eda11f1 : _GEN_736; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_738 = 11'h2e2 == io_cosIndex[10:0] ? 30'h3ed95beb : _GEN_737; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_739 = 11'h2e3 == io_cosIndex[10:0] ? 30'h3ed8a5c3 : _GEN_738; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_740 = 11'h2e4 == io_cosIndex[10:0] ? 30'h3ed7ef7a : _GEN_739; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_741 = 11'h2e5 == io_cosIndex[10:0] ? 30'h3ed73910 : _GEN_740; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_742 = 11'h2e6 == io_cosIndex[10:0] ? 30'h3ed68285 : _GEN_741; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_743 = 11'h2e7 == io_cosIndex[10:0] ? 30'h3ed5cbd8 : _GEN_742; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_744 = 11'h2e8 == io_cosIndex[10:0] ? 30'h3ed5150b : _GEN_743; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_745 = 11'h2e9 == io_cosIndex[10:0] ? 30'h3ed45e1c : _GEN_744; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_746 = 11'h2ea == io_cosIndex[10:0] ? 30'h3ed3a70d : _GEN_745; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_747 = 11'h2eb == io_cosIndex[10:0] ? 30'h3ed2efdd : _GEN_746; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_748 = 11'h2ec == io_cosIndex[10:0] ? 30'h3ed2388d : _GEN_747; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_749 = 11'h2ed == io_cosIndex[10:0] ? 30'h3ed1811c : _GEN_748; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_750 = 11'h2ee == io_cosIndex[10:0] ? 30'h3ed0c98b : _GEN_749; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_751 = 11'h2ef == io_cosIndex[10:0] ? 30'h3ed011da : _GEN_750; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_752 = 11'h2f0 == io_cosIndex[10:0] ? 30'h3ecf5a08 : _GEN_751; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_753 = 11'h2f1 == io_cosIndex[10:0] ? 30'h3ecea217 : _GEN_752; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_754 = 11'h2f2 == io_cosIndex[10:0] ? 30'h3ecdea06 : _GEN_753; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_755 = 11'h2f3 == io_cosIndex[10:0] ? 30'h3ecd31d4 : _GEN_754; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_756 = 11'h2f4 == io_cosIndex[10:0] ? 30'h3ecc7984 : _GEN_755; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_757 = 11'h2f5 == io_cosIndex[10:0] ? 30'h3ecbc113 : _GEN_756; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_758 = 11'h2f6 == io_cosIndex[10:0] ? 30'h3ecb0884 : _GEN_757; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_759 = 11'h2f7 == io_cosIndex[10:0] ? 30'h3eca4fd5 : _GEN_758; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_760 = 11'h2f8 == io_cosIndex[10:0] ? 30'h3ec99706 : _GEN_759; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_761 = 11'h2f9 == io_cosIndex[10:0] ? 30'h3ec8de19 : _GEN_760; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_762 = 11'h2fa == io_cosIndex[10:0] ? 30'h3ec8250d : _GEN_761; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_763 = 11'h2fb == io_cosIndex[10:0] ? 30'h3ec76be2 : _GEN_762; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_764 = 11'h2fc == io_cosIndex[10:0] ? 30'h3ec6b298 : _GEN_763; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_765 = 11'h2fd == io_cosIndex[10:0] ? 30'h3ec5f92f : _GEN_764; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_766 = 11'h2fe == io_cosIndex[10:0] ? 30'h3ec53fa8 : _GEN_765; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_767 = 11'h2ff == io_cosIndex[10:0] ? 30'h3ec48602 : _GEN_766; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_768 = 11'h300 == io_cosIndex[10:0] ? 30'h3ec3cc3e : _GEN_767; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_769 = 11'h301 == io_cosIndex[10:0] ? 30'h3ec3125c : _GEN_768; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_770 = 11'h302 == io_cosIndex[10:0] ? 30'h3ec2585c : _GEN_769; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_771 = 11'h303 == io_cosIndex[10:0] ? 30'h3ec19e3e : _GEN_770; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_772 = 11'h304 == io_cosIndex[10:0] ? 30'h3ec0e401 : _GEN_771; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_773 = 11'h305 == io_cosIndex[10:0] ? 30'h3ec029a8 : _GEN_772; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_774 = 11'h306 == io_cosIndex[10:0] ? 30'h3ebf6f30 : _GEN_773; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_775 = 11'h307 == io_cosIndex[10:0] ? 30'h3ebeb49b : _GEN_774; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_776 = 11'h308 == io_cosIndex[10:0] ? 30'h3ebdf9e8 : _GEN_775; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_777 = 11'h309 == io_cosIndex[10:0] ? 30'h3ebd3f19 : _GEN_776; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_778 = 11'h30a == io_cosIndex[10:0] ? 30'h3ebc842c : _GEN_777; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_779 = 11'h30b == io_cosIndex[10:0] ? 30'h3ebbc922 : _GEN_778; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_780 = 11'h30c == io_cosIndex[10:0] ? 30'h3ebb0dfb : _GEN_779; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_781 = 11'h30d == io_cosIndex[10:0] ? 30'h3eba52b7 : _GEN_780; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_782 = 11'h30e == io_cosIndex[10:0] ? 30'h3eb99756 : _GEN_781; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_783 = 11'h30f == io_cosIndex[10:0] ? 30'h3eb8dbd9 : _GEN_782; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_784 = 11'h310 == io_cosIndex[10:0] ? 30'h3eb8203f : _GEN_783; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_785 = 11'h311 == io_cosIndex[10:0] ? 30'h3eb76489 : _GEN_784; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_786 = 11'h312 == io_cosIndex[10:0] ? 30'h3eb6a8b6 : _GEN_785; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_787 = 11'h313 == io_cosIndex[10:0] ? 30'h3eb5ecc7 : _GEN_786; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_788 = 11'h314 == io_cosIndex[10:0] ? 30'h3eb530bd : _GEN_787; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_789 = 11'h315 == io_cosIndex[10:0] ? 30'h3eb47496 : _GEN_788; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_790 = 11'h316 == io_cosIndex[10:0] ? 30'h3eb3b853 : _GEN_789; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_791 = 11'h317 == io_cosIndex[10:0] ? 30'h3eb2fbf5 : _GEN_790; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_792 = 11'h318 == io_cosIndex[10:0] ? 30'h3eb23f7b : _GEN_791; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_793 = 11'h319 == io_cosIndex[10:0] ? 30'h3eb182e6 : _GEN_792; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_794 = 11'h31a == io_cosIndex[10:0] ? 30'h3eb0c635 : _GEN_793; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_795 = 11'h31b == io_cosIndex[10:0] ? 30'h3eb00969 : _GEN_794; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_796 = 11'h31c == io_cosIndex[10:0] ? 30'h3eaf4c82 : _GEN_795; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_797 = 11'h31d == io_cosIndex[10:0] ? 30'h3eae8f7f : _GEN_796; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_798 = 11'h31e == io_cosIndex[10:0] ? 30'h3eadd262 : _GEN_797; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_799 = 11'h31f == io_cosIndex[10:0] ? 30'h3ead152a : _GEN_798; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_800 = 11'h320 == io_cosIndex[10:0] ? 30'h3eac57d7 : _GEN_799; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_801 = 11'h321 == io_cosIndex[10:0] ? 30'h3eab9a6a : _GEN_800; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_802 = 11'h322 == io_cosIndex[10:0] ? 30'h3eaadce2 : _GEN_801; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_803 = 11'h323 == io_cosIndex[10:0] ? 30'h3eaa1f40 : _GEN_802; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_804 = 11'h324 == io_cosIndex[10:0] ? 30'h3ea96184 : _GEN_803; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_805 = 11'h325 == io_cosIndex[10:0] ? 30'h3ea8a3ad : _GEN_804; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_806 = 11'h326 == io_cosIndex[10:0] ? 30'h3ea7e5bd : _GEN_805; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_807 = 11'h327 == io_cosIndex[10:0] ? 30'h3ea727b2 : _GEN_806; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_808 = 11'h328 == io_cosIndex[10:0] ? 30'h3ea6698e : _GEN_807; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_809 = 11'h329 == io_cosIndex[10:0] ? 30'h3ea5ab50 : _GEN_808; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_810 = 11'h32a == io_cosIndex[10:0] ? 30'h3ea4ecf8 : _GEN_809; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_811 = 11'h32b == io_cosIndex[10:0] ? 30'h3ea42e88 : _GEN_810; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_812 = 11'h32c == io_cosIndex[10:0] ? 30'h3ea36ffd : _GEN_811; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_813 = 11'h32d == io_cosIndex[10:0] ? 30'h3ea2b15a : _GEN_812; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_814 = 11'h32e == io_cosIndex[10:0] ? 30'h3ea1f29d : _GEN_813; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_815 = 11'h32f == io_cosIndex[10:0] ? 30'h3ea133c8 : _GEN_814; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_816 = 11'h330 == io_cosIndex[10:0] ? 30'h3ea074d9 : _GEN_815; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_817 = 11'h331 == io_cosIndex[10:0] ? 30'h3e9fb5d2 : _GEN_816; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_818 = 11'h332 == io_cosIndex[10:0] ? 30'h3e9ef6b2 : _GEN_817; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_819 = 11'h333 == io_cosIndex[10:0] ? 30'h3e9e377a : _GEN_818; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_820 = 11'h334 == io_cosIndex[10:0] ? 30'h3e9d7829 : _GEN_819; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_821 = 11'h335 == io_cosIndex[10:0] ? 30'h3e9cb8c0 : _GEN_820; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_822 = 11'h336 == io_cosIndex[10:0] ? 30'h3e9bf93f : _GEN_821; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_823 = 11'h337 == io_cosIndex[10:0] ? 30'h3e9b39a5 : _GEN_822; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_824 = 11'h338 == io_cosIndex[10:0] ? 30'h3e9a79f4 : _GEN_823; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_825 = 11'h339 == io_cosIndex[10:0] ? 30'h3e99ba2b : _GEN_824; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_826 = 11'h33a == io_cosIndex[10:0] ? 30'h3e98fa4a : _GEN_825; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_827 = 11'h33b == io_cosIndex[10:0] ? 30'h3e983a52 : _GEN_826; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_828 = 11'h33c == io_cosIndex[10:0] ? 30'h3e977a42 : _GEN_827; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_829 = 11'h33d == io_cosIndex[10:0] ? 30'h3e96ba1a : _GEN_828; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_830 = 11'h33e == io_cosIndex[10:0] ? 30'h3e95f9dc : _GEN_829; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_831 = 11'h33f == io_cosIndex[10:0] ? 30'h3e953986 : _GEN_830; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_832 = 11'h340 == io_cosIndex[10:0] ? 30'h3e94791a : _GEN_831; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_833 = 11'h341 == io_cosIndex[10:0] ? 30'h3e93b896 : _GEN_832; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_834 = 11'h342 == io_cosIndex[10:0] ? 30'h3e92f7fc : _GEN_833; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_835 = 11'h343 == io_cosIndex[10:0] ? 30'h3e92374a : _GEN_834; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_836 = 11'h344 == io_cosIndex[10:0] ? 30'h3e917683 : _GEN_835; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_837 = 11'h345 == io_cosIndex[10:0] ? 30'h3e90b5a5 : _GEN_836; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_838 = 11'h346 == io_cosIndex[10:0] ? 30'h3e8ff4b0 : _GEN_837; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_839 = 11'h347 == io_cosIndex[10:0] ? 30'h3e8f33a6 : _GEN_838; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_840 = 11'h348 == io_cosIndex[10:0] ? 30'h3e8e7285 : _GEN_839; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_841 = 11'h349 == io_cosIndex[10:0] ? 30'h3e8db14e : _GEN_840; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_842 = 11'h34a == io_cosIndex[10:0] ? 30'h3e8cf002 : _GEN_841; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_843 = 11'h34b == io_cosIndex[10:0] ? 30'h3e8c2e9f : _GEN_842; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_844 = 11'h34c == io_cosIndex[10:0] ? 30'h3e8b6d28 : _GEN_843; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_845 = 11'h34d == io_cosIndex[10:0] ? 30'h3e8aab9a : _GEN_844; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_846 = 11'h34e == io_cosIndex[10:0] ? 30'h3e89e9f7 : _GEN_845; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_847 = 11'h34f == io_cosIndex[10:0] ? 30'h3e89283f : _GEN_846; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_848 = 11'h350 == io_cosIndex[10:0] ? 30'h3e886672 : _GEN_847; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_849 = 11'h351 == io_cosIndex[10:0] ? 30'h3e87a490 : _GEN_848; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_850 = 11'h352 == io_cosIndex[10:0] ? 30'h3e86e298 : _GEN_849; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_851 = 11'h353 == io_cosIndex[10:0] ? 30'h3e86208c : _GEN_850; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_852 = 11'h354 == io_cosIndex[10:0] ? 30'h3e855e6b : _GEN_851; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_853 = 11'h355 == io_cosIndex[10:0] ? 30'h3e849c36 : _GEN_852; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_854 = 11'h356 == io_cosIndex[10:0] ? 30'h3e83d9ec : _GEN_853; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_855 = 11'h357 == io_cosIndex[10:0] ? 30'h3e83178e : _GEN_854; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_856 = 11'h358 == io_cosIndex[10:0] ? 30'h3e82551c : _GEN_855; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_857 = 11'h359 == io_cosIndex[10:0] ? 30'h3e819295 : _GEN_856; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_858 = 11'h35a == io_cosIndex[10:0] ? 30'h3e80cffb : _GEN_857; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_859 = 11'h35b == io_cosIndex[10:0] ? 30'h3e800d4d : _GEN_858; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_860 = 11'h35c == io_cosIndex[10:0] ? 30'h3e7e9515 : _GEN_859; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_861 = 11'h35d == io_cosIndex[10:0] ? 30'h3e7d0f6a : _GEN_860; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_862 = 11'h35e == io_cosIndex[10:0] ? 30'h3e7b8997 : _GEN_861; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_863 = 11'h35f == io_cosIndex[10:0] ? 30'h3e7a039e : _GEN_862; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_864 = 11'h360 == io_cosIndex[10:0] ? 30'h3e787d7e : _GEN_863; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_865 = 11'h361 == io_cosIndex[10:0] ? 30'h3e76f738 : _GEN_864; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_866 = 11'h362 == io_cosIndex[10:0] ? 30'h3e7570cb : _GEN_865; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_867 = 11'h363 == io_cosIndex[10:0] ? 30'h3e73ea39 : _GEN_866; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_868 = 11'h364 == io_cosIndex[10:0] ? 30'h3e726381 : _GEN_867; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_869 = 11'h365 == io_cosIndex[10:0] ? 30'h3e70dca4 : _GEN_868; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_870 = 11'h366 == io_cosIndex[10:0] ? 30'h3e6f55a2 : _GEN_869; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_871 = 11'h367 == io_cosIndex[10:0] ? 30'h3e6dce7a : _GEN_870; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_872 = 11'h368 == io_cosIndex[10:0] ? 30'h3e6c472e : _GEN_871; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_873 = 11'h369 == io_cosIndex[10:0] ? 30'h3e6abfbe : _GEN_872; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_874 = 11'h36a == io_cosIndex[10:0] ? 30'h3e693829 : _GEN_873; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_875 = 11'h36b == io_cosIndex[10:0] ? 30'h3e67b071 : _GEN_874; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_876 = 11'h36c == io_cosIndex[10:0] ? 30'h3e662894 : _GEN_875; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_877 = 11'h36d == io_cosIndex[10:0] ? 30'h3e64a094 : _GEN_876; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_878 = 11'h36e == io_cosIndex[10:0] ? 30'h3e631871 : _GEN_877; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_879 = 11'h36f == io_cosIndex[10:0] ? 30'h3e61902b : _GEN_878; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_880 = 11'h370 == io_cosIndex[10:0] ? 30'h3e6007c2 : _GEN_879; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_881 = 11'h371 == io_cosIndex[10:0] ? 30'h3e5e7f36 : _GEN_880; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_882 = 11'h372 == io_cosIndex[10:0] ? 30'h3e5cf688 : _GEN_881; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_883 = 11'h373 == io_cosIndex[10:0] ? 30'h3e5b6db8 : _GEN_882; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_884 = 11'h374 == io_cosIndex[10:0] ? 30'h3e59e4c6 : _GEN_883; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_885 = 11'h375 == io_cosIndex[10:0] ? 30'h3e585bb3 : _GEN_884; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_886 = 11'h376 == io_cosIndex[10:0] ? 30'h3e56d27e : _GEN_885; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_887 = 11'h377 == io_cosIndex[10:0] ? 30'h3e554928 : _GEN_886; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_888 = 11'h378 == io_cosIndex[10:0] ? 30'h3e53bfb1 : _GEN_887; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_889 = 11'h379 == io_cosIndex[10:0] ? 30'h3e52361a : _GEN_888; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_890 = 11'h37a == io_cosIndex[10:0] ? 30'h3e50ac61 : _GEN_889; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_891 = 11'h37b == io_cosIndex[10:0] ? 30'h3e4f2289 : _GEN_890; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_892 = 11'h37c == io_cosIndex[10:0] ? 30'h3e4d9891 : _GEN_891; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_893 = 11'h37d == io_cosIndex[10:0] ? 30'h3e4c0e79 : _GEN_892; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_894 = 11'h37e == io_cosIndex[10:0] ? 30'h3e4a8442 : _GEN_893; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_895 = 11'h37f == io_cosIndex[10:0] ? 30'h3e48f9eb : _GEN_894; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_896 = 11'h380 == io_cosIndex[10:0] ? 30'h3e476f76 : _GEN_895; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_897 = 11'h381 == io_cosIndex[10:0] ? 30'h3e45e4e1 : _GEN_896; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_898 = 11'h382 == io_cosIndex[10:0] ? 30'h3e445a2e : _GEN_897; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_899 = 11'h383 == io_cosIndex[10:0] ? 30'h3e42cf5d : _GEN_898; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_900 = 11'h384 == io_cosIndex[10:0] ? 30'h3e41446e : _GEN_899; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_901 = 11'h385 == io_cosIndex[10:0] ? 30'h3e3fb961 : _GEN_900; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_902 = 11'h386 == io_cosIndex[10:0] ? 30'h3e3e2e36 : _GEN_901; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_903 = 11'h387 == io_cosIndex[10:0] ? 30'h3e3ca2ee : _GEN_902; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_904 = 11'h388 == io_cosIndex[10:0] ? 30'h3e3b1789 : _GEN_903; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_905 = 11'h389 == io_cosIndex[10:0] ? 30'h3e398c07 : _GEN_904; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_906 = 11'h38a == io_cosIndex[10:0] ? 30'h3e380068 : _GEN_905; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_907 = 11'h38b == io_cosIndex[10:0] ? 30'h3e3674ad : _GEN_906; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_908 = 11'h38c == io_cosIndex[10:0] ? 30'h3e34e8d6 : _GEN_907; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_909 = 11'h38d == io_cosIndex[10:0] ? 30'h3e335ce3 : _GEN_908; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_910 = 11'h38e == io_cosIndex[10:0] ? 30'h3e31d0d4 : _GEN_909; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_911 = 11'h38f == io_cosIndex[10:0] ? 30'h3e3044aa : _GEN_910; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_912 = 11'h390 == io_cosIndex[10:0] ? 30'h3e2eb864 : _GEN_911; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_913 = 11'h391 == io_cosIndex[10:0] ? 30'h3e2d2c04 : _GEN_912; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_914 = 11'h392 == io_cosIndex[10:0] ? 30'h3e2b9f89 : _GEN_913; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_915 = 11'h393 == io_cosIndex[10:0] ? 30'h3e2a12f3 : _GEN_914; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_916 = 11'h394 == io_cosIndex[10:0] ? 30'h3e288644 : _GEN_915; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_917 = 11'h395 == io_cosIndex[10:0] ? 30'h3e26f97a : _GEN_916; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_918 = 11'h396 == io_cosIndex[10:0] ? 30'h3e256c96 : _GEN_917; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_919 = 11'h397 == io_cosIndex[10:0] ? 30'h3e23df99 : _GEN_918; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_920 = 11'h398 == io_cosIndex[10:0] ? 30'h3e225283 : _GEN_919; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_921 = 11'h399 == io_cosIndex[10:0] ? 30'h3e20c553 : _GEN_920; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_922 = 11'h39a == io_cosIndex[10:0] ? 30'h3e1f380b : _GEN_921; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_923 = 11'h39b == io_cosIndex[10:0] ? 30'h3e1daaaa : _GEN_922; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_924 = 11'h39c == io_cosIndex[10:0] ? 30'h3e1c1d31 : _GEN_923; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_925 = 11'h39d == io_cosIndex[10:0] ? 30'h3e1a8fa0 : _GEN_924; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_926 = 11'h39e == io_cosIndex[10:0] ? 30'h3e1901f7 : _GEN_925; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_927 = 11'h39f == io_cosIndex[10:0] ? 30'h3e177436 : _GEN_926; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_928 = 11'h3a0 == io_cosIndex[10:0] ? 30'h3e15e65e : _GEN_927; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_929 = 11'h3a1 == io_cosIndex[10:0] ? 30'h3e14586f : _GEN_928; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_930 = 11'h3a2 == io_cosIndex[10:0] ? 30'h3e12ca69 : _GEN_929; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_931 = 11'h3a3 == io_cosIndex[10:0] ? 30'h3e113c4d : _GEN_930; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_932 = 11'h3a4 == io_cosIndex[10:0] ? 30'h3e0fae1a : _GEN_931; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_933 = 11'h3a5 == io_cosIndex[10:0] ? 30'h3e0e1fd0 : _GEN_932; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_934 = 11'h3a6 == io_cosIndex[10:0] ? 30'h3e0c9171 : _GEN_933; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_935 = 11'h3a7 == io_cosIndex[10:0] ? 30'h3e0b02fc : _GEN_934; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_936 = 11'h3a8 == io_cosIndex[10:0] ? 30'h3e097472 : _GEN_935; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_937 = 11'h3a9 == io_cosIndex[10:0] ? 30'h3e07e5d2 : _GEN_936; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_938 = 11'h3aa == io_cosIndex[10:0] ? 30'h3e06571e : _GEN_937; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_939 = 11'h3ab == io_cosIndex[10:0] ? 30'h3e04c855 : _GEN_938; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_940 = 11'h3ac == io_cosIndex[10:0] ? 30'h3e033977 : _GEN_939; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_941 = 11'h3ad == io_cosIndex[10:0] ? 30'h3e01aa85 : _GEN_940; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_942 = 11'h3ae == io_cosIndex[10:0] ? 30'h3e001b7f : _GEN_941; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_943 = 11'h3af == io_cosIndex[10:0] ? 30'h3dfd18cb : _GEN_942; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_944 = 11'h3b0 == io_cosIndex[10:0] ? 30'h3df9fa70 : _GEN_943; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_945 = 11'h3b1 == io_cosIndex[10:0] ? 30'h3df6dbef : _GEN_944; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_946 = 11'h3b2 == io_cosIndex[10:0] ? 30'h3df3bd48 : _GEN_945; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_947 = 11'h3b3 == io_cosIndex[10:0] ? 30'h3df09e7b : _GEN_946; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_948 = 11'h3b4 == io_cosIndex[10:0] ? 30'h3ded7f8a : _GEN_947; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_949 = 11'h3b5 == io_cosIndex[10:0] ? 30'h3dea6073 : _GEN_948; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_950 = 11'h3b6 == io_cosIndex[10:0] ? 30'h3de74138 : _GEN_949; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_951 = 11'h3b7 == io_cosIndex[10:0] ? 30'h3de421da : _GEN_950; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_952 = 11'h3b8 == io_cosIndex[10:0] ? 30'h3de10259 : _GEN_951; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_953 = 11'h3b9 == io_cosIndex[10:0] ? 30'h3ddde2b4 : _GEN_952; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_954 = 11'h3ba == io_cosIndex[10:0] ? 30'h3ddac2ee : _GEN_953; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_955 = 11'h3bb == io_cosIndex[10:0] ? 30'h3dd7a305 : _GEN_954; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_956 = 11'h3bc == io_cosIndex[10:0] ? 30'h3dd482fc : _GEN_955; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_957 = 11'h3bd == io_cosIndex[10:0] ? 30'h3dd162d2 : _GEN_956; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_958 = 11'h3be == io_cosIndex[10:0] ? 30'h3dce4287 : _GEN_957; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_959 = 11'h3bf == io_cosIndex[10:0] ? 30'h3dcb221d : _GEN_958; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_960 = 11'h3c0 == io_cosIndex[10:0] ? 30'h3dc80193 : _GEN_959; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_961 = 11'h3c1 == io_cosIndex[10:0] ? 30'h3dc4e0ea : _GEN_960; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_962 = 11'h3c2 == io_cosIndex[10:0] ? 30'h3dc1c023 : _GEN_961; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_963 = 11'h3c3 == io_cosIndex[10:0] ? 30'h3dbe9f3e : _GEN_962; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_964 = 11'h3c4 == io_cosIndex[10:0] ? 30'h3dbb7e3c : _GEN_963; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_965 = 11'h3c5 == io_cosIndex[10:0] ? 30'h3db85d1d : _GEN_964; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_966 = 11'h3c6 == io_cosIndex[10:0] ? 30'h3db53be1 : _GEN_965; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_967 = 11'h3c7 == io_cosIndex[10:0] ? 30'h3db21a89 : _GEN_966; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_968 = 11'h3c8 == io_cosIndex[10:0] ? 30'h3daef916 : _GEN_967; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_969 = 11'h3c9 == io_cosIndex[10:0] ? 30'h3dabd788 : _GEN_968; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_970 = 11'h3ca == io_cosIndex[10:0] ? 30'h3da8b5df : _GEN_969; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_971 = 11'h3cb == io_cosIndex[10:0] ? 30'h3da5941d : _GEN_970; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_972 = 11'h3cc == io_cosIndex[10:0] ? 30'h3da27240 : _GEN_971; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_973 = 11'h3cd == io_cosIndex[10:0] ? 30'h3d9f504b : _GEN_972; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_974 = 11'h3ce == io_cosIndex[10:0] ? 30'h3d9c2e3d : _GEN_973; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_975 = 11'h3cf == io_cosIndex[10:0] ? 30'h3d990c17 : _GEN_974; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_976 = 11'h3d0 == io_cosIndex[10:0] ? 30'h3d95e9da : _GEN_975; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_977 = 11'h3d1 == io_cosIndex[10:0] ? 30'h3d92c785 : _GEN_976; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_978 = 11'h3d2 == io_cosIndex[10:0] ? 30'h3d8fa51a : _GEN_977; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_979 = 11'h3d3 == io_cosIndex[10:0] ? 30'h3d8c8298 : _GEN_978; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_980 = 11'h3d4 == io_cosIndex[10:0] ? 30'h3d896001 : _GEN_979; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_981 = 11'h3d5 == io_cosIndex[10:0] ? 30'h3d863d55 : _GEN_980; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_982 = 11'h3d6 == io_cosIndex[10:0] ? 30'h3d831a94 : _GEN_981; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_983 = 11'h3d7 == io_cosIndex[10:0] ? 30'h3d7fef7c : _GEN_982; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_984 = 11'h3d8 == io_cosIndex[10:0] ? 30'h3d79a9aa : _GEN_983; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_985 = 11'h3d9 == io_cosIndex[10:0] ? 30'h3d7363b2 : _GEN_984; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_986 = 11'h3da == io_cosIndex[10:0] ? 30'h3d6d1d93 : _GEN_985; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_987 = 11'h3db == io_cosIndex[10:0] ? 30'h3d66d751 : _GEN_986; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_988 = 11'h3dc == io_cosIndex[10:0] ? 30'h3d6090ea : _GEN_987; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_989 = 11'h3dd == io_cosIndex[10:0] ? 30'h3d5a4a61 : _GEN_988; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_990 = 11'h3de == io_cosIndex[10:0] ? 30'h3d5403b6 : _GEN_989; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_991 = 11'h3df == io_cosIndex[10:0] ? 30'h3d4dbceb : _GEN_990; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_992 = 11'h3e0 == io_cosIndex[10:0] ? 30'h3d477600 : _GEN_991; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_993 = 11'h3e1 == io_cosIndex[10:0] ? 30'h3d412ef6 : _GEN_992; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_994 = 11'h3e2 == io_cosIndex[10:0] ? 30'h3d3ae7ce : _GEN_993; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_995 = 11'h3e3 == io_cosIndex[10:0] ? 30'h3d34a089 : _GEN_994; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_996 = 11'h3e4 == io_cosIndex[10:0] ? 30'h3d2e5929 : _GEN_995; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_997 = 11'h3e5 == io_cosIndex[10:0] ? 30'h3d2811ad : _GEN_996; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_998 = 11'h3e6 == io_cosIndex[10:0] ? 30'h3d21ca18 : _GEN_997; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_999 = 11'h3e7 == io_cosIndex[10:0] ? 30'h3d1b826a : _GEN_998; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1000 = 11'h3e8 == io_cosIndex[10:0] ? 30'h3d153aa4 : _GEN_999; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1001 = 11'h3e9 == io_cosIndex[10:0] ? 30'h3d0ef2c6 : _GEN_1000; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1002 = 11'h3ea == io_cosIndex[10:0] ? 30'h3d08aad3 : _GEN_1001; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1003 = 11'h3eb == io_cosIndex[10:0] ? 30'h3d0262cb : _GEN_1002; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1004 = 11'h3ec == io_cosIndex[10:0] ? 30'h3cf8355c : _GEN_1003; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1005 = 11'h3ed == io_cosIndex[10:0] ? 30'h3ceba4fd : _GEN_1004; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1006 = 11'h3ee == io_cosIndex[10:0] ? 30'h3cdf1479 : _GEN_1005; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1007 = 11'h3ef == io_cosIndex[10:0] ? 30'h3cd283d3 : _GEN_1006; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1008 = 11'h3f0 == io_cosIndex[10:0] ? 30'h3cc5f30c : _GEN_1007; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1009 = 11'h3f1 == io_cosIndex[10:0] ? 30'h3cb96227 : _GEN_1008; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1010 = 11'h3f2 == io_cosIndex[10:0] ? 30'h3cacd125 : _GEN_1009; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1011 = 11'h3f3 == io_cosIndex[10:0] ? 30'h3ca04008 : _GEN_1010; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1012 = 11'h3f4 == io_cosIndex[10:0] ? 30'h3c93aed3 : _GEN_1011; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1013 = 11'h3f5 == io_cosIndex[10:0] ? 30'h3c871d87 : _GEN_1012; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1014 = 11'h3f6 == io_cosIndex[10:0] ? 30'h3c75184d : _GEN_1013; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1015 = 11'h3f7 == io_cosIndex[10:0] ? 30'h3c5bf566 : _GEN_1014; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1016 = 11'h3f8 == io_cosIndex[10:0] ? 30'h3c42d25c : _GEN_1015; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1017 = 11'h3f9 == io_cosIndex[10:0] ? 30'h3c29af35 : _GEN_1016; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1018 = 11'h3fa == io_cosIndex[10:0] ? 30'h3c108bf3 : _GEN_1017; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1019 = 11'h3fb == io_cosIndex[10:0] ? 30'h3beed136 : _GEN_1018; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1020 = 11'h3fc == io_cosIndex[10:0] ? 30'h3bbc8a61 : _GEN_1019; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1021 = 11'h3fd == io_cosIndex[10:0] ? 30'h3b8a4370 : _GEN_1020; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1022 = 11'h3fe == io_cosIndex[10:0] ? 30'h3b2ff8d1 : _GEN_1021; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1023 = 11'h3ff == io_cosIndex[10:0] ? 30'h3a96d54f : _GEN_1022; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1024 = 11'h400 == io_cosIndex[10:0] ? 30'h0 : _GEN_1023; // @[LUTbank.scala 293:{21,21}]
  wire [29:0] _GEN_1026 = 11'h1 == io_sinIndex[10:0] ? 30'h3ac91c67 : 30'h0; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1027 = 11'h2 == io_sinIndex[10:0] ? 30'h3b491c58 : _GEN_1026; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1028 = 11'h3 == io_sinIndex[10:0] ? 30'h3b96d52e : _GEN_1027; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1029 = 11'h4 == io_sinIndex[10:0] ? 30'h3bc91c1a : _GEN_1028; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1030 = 11'h5 == io_sinIndex[10:0] ? 30'h3bfb62e6 : _GEN_1029; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1031 = 11'h6 == io_sinIndex[10:0] ? 30'h3c16d4c6 : _GEN_1030; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1032 = 11'h7 == io_sinIndex[10:0] ? 30'h3c2ff801 : _GEN_1031; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1033 = 11'h8 == io_sinIndex[10:0] ? 30'h3c491b21 : _GEN_1032; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1034 = 11'h9 == io_sinIndex[10:0] ? 30'h3c623e23 : _GEN_1033; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1035 = 11'ha == io_sinIndex[10:0] ? 30'h3c7b6101 : _GEN_1034; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1036 = 11'hb == io_sinIndex[10:0] ? 30'h3c8a41dc : _GEN_1035; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1037 = 11'hc == io_sinIndex[10:0] ? 30'h3c96d323 : _GEN_1036; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1038 = 11'hd == io_sinIndex[10:0] ? 30'h3ca36452 : _GEN_1037; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1039 = 11'he == io_sinIndex[10:0] ? 30'h3caff568 : _GEN_1038; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1040 = 11'hf == io_sinIndex[10:0] ? 30'h3cbc8663 : _GEN_1039; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1041 = 11'h10 == io_sinIndex[10:0] ? 30'h3cc91741 : _GEN_1040; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1042 = 11'h11 == io_sinIndex[10:0] ? 30'h3cd5a7ff : _GEN_1041; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1043 = 11'h12 == io_sinIndex[10:0] ? 30'h3ce2389d : _GEN_1042; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1044 = 11'h13 == io_sinIndex[10:0] ? 30'h3ceec918 : _GEN_1043; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1045 = 11'h14 == io_sinIndex[10:0] ? 30'h3cfb596e : _GEN_1044; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1046 = 11'h15 == io_sinIndex[10:0] ? 30'h3d03f4cf : _GEN_1045; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1047 = 11'h16 == io_sinIndex[10:0] ? 30'h3d0a3cd2 : _GEN_1046; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1048 = 11'h17 == io_sinIndex[10:0] ? 30'h3d1084c0 : _GEN_1047; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1049 = 11'h18 == io_sinIndex[10:0] ? 30'h3d16cc97 : _GEN_1048; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1050 = 11'h19 == io_sinIndex[10:0] ? 30'h3d1d1458 : _GEN_1049; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1051 = 11'h1a == io_sinIndex[10:0] ? 30'h3d235c00 : _GEN_1050; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1052 = 11'h1b == io_sinIndex[10:0] ? 30'h3d29a38f : _GEN_1051; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1053 = 11'h1c == io_sinIndex[10:0] ? 30'h3d2feb04 : _GEN_1052; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1054 = 11'h1d == io_sinIndex[10:0] ? 30'h3d36325d : _GEN_1053; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1055 = 11'h1e == io_sinIndex[10:0] ? 30'h3d3c799b : _GEN_1054; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1056 = 11'h1f == io_sinIndex[10:0] ? 30'h3d42c0bb : _GEN_1055; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1057 = 11'h20 == io_sinIndex[10:0] ? 30'h3d4907bd : _GEN_1056; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1058 = 11'h21 == io_sinIndex[10:0] ? 30'h3d4f4ea1 : _GEN_1057; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1059 = 11'h22 == io_sinIndex[10:0] ? 30'h3d559564 : _GEN_1058; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1060 = 11'h23 == io_sinIndex[10:0] ? 30'h3d5bdc07 : _GEN_1059; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1061 = 11'h24 == io_sinIndex[10:0] ? 30'h3d622287 : _GEN_1060; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1062 = 11'h25 == io_sinIndex[10:0] ? 30'h3d6868e5 : _GEN_1061; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1063 = 11'h26 == io_sinIndex[10:0] ? 30'h3d6eaf1e : _GEN_1062; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1064 = 11'h27 == io_sinIndex[10:0] ? 30'h3d74f533 : _GEN_1063; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1065 = 11'h28 == io_sinIndex[10:0] ? 30'h3d7b3b22 : _GEN_1064; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1066 = 11'h29 == io_sinIndex[10:0] ? 30'h3d80c075 : _GEN_1065; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1067 = 11'h2a == io_sinIndex[10:0] ? 30'h3d83e346 : _GEN_1066; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1068 = 11'h2b == io_sinIndex[10:0] ? 30'h3d870602 : _GEN_1067; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1069 = 11'h2c == io_sinIndex[10:0] ? 30'h3d8a28a9 : _GEN_1068; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1070 = 11'h2d == io_sinIndex[10:0] ? 30'h3d8d4b3b : _GEN_1069; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1071 = 11'h2e == io_sinIndex[10:0] ? 30'h3d906db7 : _GEN_1070; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1072 = 11'h2f == io_sinIndex[10:0] ? 30'h3d93901c : _GEN_1071; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1073 = 11'h30 == io_sinIndex[10:0] ? 30'h3d96b26b : _GEN_1072; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1074 = 11'h31 == io_sinIndex[10:0] ? 30'h3d99d4a3 : _GEN_1073; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1075 = 11'h32 == io_sinIndex[10:0] ? 30'h3d9cf6c3 : _GEN_1074; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1076 = 11'h33 == io_sinIndex[10:0] ? 30'h3da018cb : _GEN_1075; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1077 = 11'h34 == io_sinIndex[10:0] ? 30'h3da33aba : _GEN_1076; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1078 = 11'h35 == io_sinIndex[10:0] ? 30'h3da65c90 : _GEN_1077; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1079 = 11'h36 == io_sinIndex[10:0] ? 30'h3da97e4c : _GEN_1078; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1080 = 11'h37 == io_sinIndex[10:0] ? 30'h3dac9fee : _GEN_1079; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1081 = 11'h38 == io_sinIndex[10:0] ? 30'h3dafc176 : _GEN_1080; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1082 = 11'h39 == io_sinIndex[10:0] ? 30'h3db2e2e2 : _GEN_1081; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1083 = 11'h3a == io_sinIndex[10:0] ? 30'h3db60433 : _GEN_1082; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1084 = 11'h3b == io_sinIndex[10:0] ? 30'h3db92567 : _GEN_1083; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1085 = 11'h3c == io_sinIndex[10:0] ? 30'h3dbc467f : _GEN_1084; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1086 = 11'h3d == io_sinIndex[10:0] ? 30'h3dbf677a : _GEN_1085; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1087 = 11'h3e == io_sinIndex[10:0] ? 30'h3dc28858 : _GEN_1086; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1088 = 11'h3f == io_sinIndex[10:0] ? 30'h3dc5a917 : _GEN_1087; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1089 = 11'h40 == io_sinIndex[10:0] ? 30'h3dc8c9b8 : _GEN_1088; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1090 = 11'h41 == io_sinIndex[10:0] ? 30'h3dcbea3a : _GEN_1089; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1091 = 11'h42 == io_sinIndex[10:0] ? 30'h3dcf0a9d : _GEN_1090; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1092 = 11'h43 == io_sinIndex[10:0] ? 30'h3dd22adf : _GEN_1091; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1093 = 11'h44 == io_sinIndex[10:0] ? 30'h3dd54b01 : _GEN_1092; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1094 = 11'h45 == io_sinIndex[10:0] ? 30'h3dd86b03 : _GEN_1093; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1095 = 11'h46 == io_sinIndex[10:0] ? 30'h3ddb8ae3 : _GEN_1094; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1096 = 11'h47 == io_sinIndex[10:0] ? 30'h3ddeaaa1 : _GEN_1095; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1097 = 11'h48 == io_sinIndex[10:0] ? 30'h3de1ca3c : _GEN_1096; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1098 = 11'h49 == io_sinIndex[10:0] ? 30'h3de4e9b5 : _GEN_1097; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1099 = 11'h4a == io_sinIndex[10:0] ? 30'h3de8090a : _GEN_1098; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1100 = 11'h4b == io_sinIndex[10:0] ? 30'h3deb283c : _GEN_1099; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1101 = 11'h4c == io_sinIndex[10:0] ? 30'h3dee474a : _GEN_1100; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1102 = 11'h4d == io_sinIndex[10:0] ? 30'h3df16632 : _GEN_1101; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1103 = 11'h4e == io_sinIndex[10:0] ? 30'h3df484f6 : _GEN_1102; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1104 = 11'h4f == io_sinIndex[10:0] ? 30'h3df7a393 : _GEN_1103; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1105 = 11'h50 == io_sinIndex[10:0] ? 30'h3dfac20b : _GEN_1104; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1106 = 11'h51 == io_sinIndex[10:0] ? 30'h3dfde05b : _GEN_1105; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1107 = 11'h52 == io_sinIndex[10:0] ? 30'h3e007f43 : _GEN_1106; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1108 = 11'h53 == io_sinIndex[10:0] ? 30'h3e020e43 : _GEN_1107; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1109 = 11'h54 == io_sinIndex[10:0] ? 30'h3e039d30 : _GEN_1108; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1110 = 11'h55 == io_sinIndex[10:0] ? 30'h3e052c09 : _GEN_1109; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1111 = 11'h56 == io_sinIndex[10:0] ? 30'h3e06bacd : _GEN_1110; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1112 = 11'h57 == io_sinIndex[10:0] ? 30'h3e08497c : _GEN_1111; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1113 = 11'h58 == io_sinIndex[10:0] ? 30'h3e09d817 : _GEN_1112; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1114 = 11'h59 == io_sinIndex[10:0] ? 30'h3e0b669c : _GEN_1113; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1115 = 11'h5a == io_sinIndex[10:0] ? 30'h3e0cf50b : _GEN_1114; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1116 = 11'h5b == io_sinIndex[10:0] ? 30'h3e0e8365 : _GEN_1115; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1117 = 11'h5c == io_sinIndex[10:0] ? 30'h3e1011a8 : _GEN_1116; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1118 = 11'h5d == io_sinIndex[10:0] ? 30'h3e119fd6 : _GEN_1117; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1119 = 11'h5e == io_sinIndex[10:0] ? 30'h3e132ded : _GEN_1118; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1120 = 11'h5f == io_sinIndex[10:0] ? 30'h3e14bbed : _GEN_1119; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1121 = 11'h60 == io_sinIndex[10:0] ? 30'h3e1649d7 : _GEN_1120; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1122 = 11'h61 == io_sinIndex[10:0] ? 30'h3e17d7a9 : _GEN_1121; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1123 = 11'h62 == io_sinIndex[10:0] ? 30'h3e196564 : _GEN_1122; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1124 = 11'h63 == io_sinIndex[10:0] ? 30'h3e1af307 : _GEN_1123; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1125 = 11'h64 == io_sinIndex[10:0] ? 30'h3e1c8092 : _GEN_1124; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1126 = 11'h65 == io_sinIndex[10:0] ? 30'h3e1e0e05 : _GEN_1125; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1127 = 11'h66 == io_sinIndex[10:0] ? 30'h3e1f9b60 : _GEN_1126; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1128 = 11'h67 == io_sinIndex[10:0] ? 30'h3e2128a2 : _GEN_1127; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1129 = 11'h68 == io_sinIndex[10:0] ? 30'h3e22b5cb : _GEN_1128; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1130 = 11'h69 == io_sinIndex[10:0] ? 30'h3e2442db : _GEN_1129; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1131 = 11'h6a == io_sinIndex[10:0] ? 30'h3e25cfd2 : _GEN_1130; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1132 = 11'h6b == io_sinIndex[10:0] ? 30'h3e275caf : _GEN_1131; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1133 = 11'h6c == io_sinIndex[10:0] ? 30'h3e28e972 : _GEN_1132; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1134 = 11'h6d == io_sinIndex[10:0] ? 30'h3e2a761b : _GEN_1133; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1135 = 11'h6e == io_sinIndex[10:0] ? 30'h3e2c02aa : _GEN_1134; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1136 = 11'h6f == io_sinIndex[10:0] ? 30'h3e2d8f1f : _GEN_1135; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1137 = 11'h70 == io_sinIndex[10:0] ? 30'h3e2f1b78 : _GEN_1136; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1138 = 11'h71 == io_sinIndex[10:0] ? 30'h3e30a7b7 : _GEN_1137; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1139 = 11'h72 == io_sinIndex[10:0] ? 30'h3e3233da : _GEN_1138; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1140 = 11'h73 == io_sinIndex[10:0] ? 30'h3e33bfe2 : _GEN_1139; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1141 = 11'h74 == io_sinIndex[10:0] ? 30'h3e354bce : _GEN_1140; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1142 = 11'h75 == io_sinIndex[10:0] ? 30'h3e36d79e : _GEN_1141; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1143 = 11'h76 == io_sinIndex[10:0] ? 30'h3e386352 : _GEN_1142; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1144 = 11'h77 == io_sinIndex[10:0] ? 30'h3e39eeea : _GEN_1143; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1145 = 11'h78 == io_sinIndex[10:0] ? 30'h3e3b7a65 : _GEN_1144; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1146 = 11'h79 == io_sinIndex[10:0] ? 30'h3e3d05c3 : _GEN_1145; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1147 = 11'h7a == io_sinIndex[10:0] ? 30'h3e3e9103 : _GEN_1146; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1148 = 11'h7b == io_sinIndex[10:0] ? 30'h3e401c27 : _GEN_1147; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1149 = 11'h7c == io_sinIndex[10:0] ? 30'h3e41a72c : _GEN_1148; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1150 = 11'h7d == io_sinIndex[10:0] ? 30'h3e433214 : _GEN_1149; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1151 = 11'h7e == io_sinIndex[10:0] ? 30'h3e44bcde : _GEN_1150; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1152 = 11'h7f == io_sinIndex[10:0] ? 30'h3e464789 : _GEN_1151; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1153 = 11'h80 == io_sinIndex[10:0] ? 30'h3e47d216 : _GEN_1152; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1154 = 11'h81 == io_sinIndex[10:0] ? 30'h3e495c84 : _GEN_1153; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1155 = 11'h82 == io_sinIndex[10:0] ? 30'h3e4ae6d3 : _GEN_1154; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1156 = 11'h83 == io_sinIndex[10:0] ? 30'h3e4c7102 : _GEN_1155; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1157 = 11'h84 == io_sinIndex[10:0] ? 30'h3e4dfb12 : _GEN_1156; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1158 = 11'h85 == io_sinIndex[10:0] ? 30'h3e4f8502 : _GEN_1157; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1159 = 11'h86 == io_sinIndex[10:0] ? 30'h3e510ed3 : _GEN_1158; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1160 = 11'h87 == io_sinIndex[10:0] ? 30'h3e529882 : _GEN_1159; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1161 = 11'h88 == io_sinIndex[10:0] ? 30'h3e542212 : _GEN_1160; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1162 = 11'h89 == io_sinIndex[10:0] ? 30'h3e55ab81 : _GEN_1161; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1163 = 11'h8a == io_sinIndex[10:0] ? 30'h3e5734ce : _GEN_1162; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1164 = 11'h8b == io_sinIndex[10:0] ? 30'h3e58bdfb : _GEN_1163; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1165 = 11'h8c == io_sinIndex[10:0] ? 30'h3e5a4706 : _GEN_1164; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1166 = 11'h8d == io_sinIndex[10:0] ? 30'h3e5bcfef : _GEN_1165; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1167 = 11'h8e == io_sinIndex[10:0] ? 30'h3e5d58b7 : _GEN_1166; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1168 = 11'h8f == io_sinIndex[10:0] ? 30'h3e5ee15c : _GEN_1167; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1169 = 11'h90 == io_sinIndex[10:0] ? 30'h3e6069df : _GEN_1168; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1170 = 11'h91 == io_sinIndex[10:0] ? 30'h3e61f240 : _GEN_1169; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1171 = 11'h92 == io_sinIndex[10:0] ? 30'h3e637a7d : _GEN_1170; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1172 = 11'h93 == io_sinIndex[10:0] ? 30'h3e650298 : _GEN_1171; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1173 = 11'h94 == io_sinIndex[10:0] ? 30'h3e668a8f : _GEN_1172; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1174 = 11'h95 == io_sinIndex[10:0] ? 30'h3e681262 : _GEN_1173; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1175 = 11'h96 == io_sinIndex[10:0] ? 30'h3e699a12 : _GEN_1174; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1176 = 11'h97 == io_sinIndex[10:0] ? 30'h3e6b219d : _GEN_1175; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1177 = 11'h98 == io_sinIndex[10:0] ? 30'h3e6ca905 : _GEN_1176; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1178 = 11'h99 == io_sinIndex[10:0] ? 30'h3e6e3048 : _GEN_1177; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1179 = 11'h9a == io_sinIndex[10:0] ? 30'h3e6fb766 : _GEN_1178; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1180 = 11'h9b == io_sinIndex[10:0] ? 30'h3e713e5f : _GEN_1179; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1181 = 11'h9c == io_sinIndex[10:0] ? 30'h3e72c533 : _GEN_1180; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1182 = 11'h9d == io_sinIndex[10:0] ? 30'h3e744be1 : _GEN_1181; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1183 = 11'h9e == io_sinIndex[10:0] ? 30'h3e75d26a : _GEN_1182; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1184 = 11'h9f == io_sinIndex[10:0] ? 30'h3e7758cd : _GEN_1183; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1185 = 11'ha0 == io_sinIndex[10:0] ? 30'h3e78df09 : _GEN_1184; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1186 = 11'ha1 == io_sinIndex[10:0] ? 30'h3e7a6520 : _GEN_1185; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1187 = 11'ha2 == io_sinIndex[10:0] ? 30'h3e7beb0f : _GEN_1186; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1188 = 11'ha3 == io_sinIndex[10:0] ? 30'h3e7d70d8 : _GEN_1187; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1189 = 11'ha4 == io_sinIndex[10:0] ? 30'h3e7ef67a : _GEN_1188; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1190 = 11'ha5 == io_sinIndex[10:0] ? 30'h3e803dfa : _GEN_1189; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1191 = 11'ha6 == io_sinIndex[10:0] ? 30'h3e8100a3 : _GEN_1190; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1192 = 11'ha7 == io_sinIndex[10:0] ? 30'h3e81c339 : _GEN_1191; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1193 = 11'ha8 == io_sinIndex[10:0] ? 30'h3e8285ba : _GEN_1192; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1194 = 11'ha9 == io_sinIndex[10:0] ? 30'h3e834828 : _GEN_1193; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1195 = 11'haa == io_sinIndex[10:0] ? 30'h3e840a81 : _GEN_1194; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1196 = 11'hab == io_sinIndex[10:0] ? 30'h3e84ccc5 : _GEN_1195; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1197 = 11'hac == io_sinIndex[10:0] ? 30'h3e858ef6 : _GEN_1196; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1198 = 11'had == io_sinIndex[10:0] ? 30'h3e865111 : _GEN_1197; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1199 = 11'hae == io_sinIndex[10:0] ? 30'h3e871318 : _GEN_1198; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1200 = 11'haf == io_sinIndex[10:0] ? 30'h3e87d50a : _GEN_1199; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1201 = 11'hb0 == io_sinIndex[10:0] ? 30'h3e8896e7 : _GEN_1200; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1202 = 11'hb1 == io_sinIndex[10:0] ? 30'h3e8958af : _GEN_1201; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1203 = 11'hb2 == io_sinIndex[10:0] ? 30'h3e8a1a62 : _GEN_1202; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1204 = 11'hb3 == io_sinIndex[10:0] ? 30'h3e8adbff : _GEN_1203; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1205 = 11'hb4 == io_sinIndex[10:0] ? 30'h3e8b9d88 : _GEN_1204; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1206 = 11'hb5 == io_sinIndex[10:0] ? 30'h3e8c5efa : _GEN_1205; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1207 = 11'hb6 == io_sinIndex[10:0] ? 30'h3e8d2057 : _GEN_1206; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1208 = 11'hb7 == io_sinIndex[10:0] ? 30'h3e8de19e : _GEN_1207; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1209 = 11'hb8 == io_sinIndex[10:0] ? 30'h3e8ea2cf : _GEN_1208; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1210 = 11'hb9 == io_sinIndex[10:0] ? 30'h3e8f63ea : _GEN_1209; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1211 = 11'hba == io_sinIndex[10:0] ? 30'h3e9024ef : _GEN_1210; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1212 = 11'hbb == io_sinIndex[10:0] ? 30'h3e90e5de : _GEN_1211; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1213 = 11'hbc == io_sinIndex[10:0] ? 30'h3e91a6b7 : _GEN_1212; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1214 = 11'hbd == io_sinIndex[10:0] ? 30'h3e926779 : _GEN_1213; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1215 = 11'hbe == io_sinIndex[10:0] ? 30'h3e932824 : _GEN_1214; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1216 = 11'hbf == io_sinIndex[10:0] ? 30'h3e93e8b9 : _GEN_1215; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1217 = 11'hc0 == io_sinIndex[10:0] ? 30'h3e94a937 : _GEN_1216; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1218 = 11'hc1 == io_sinIndex[10:0] ? 30'h3e95699e : _GEN_1217; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1219 = 11'hc2 == io_sinIndex[10:0] ? 30'h3e9629ee : _GEN_1218; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1220 = 11'hc3 == io_sinIndex[10:0] ? 30'h3e96ea26 : _GEN_1219; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1221 = 11'hc4 == io_sinIndex[10:0] ? 30'h3e97aa48 : _GEN_1220; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1222 = 11'hc5 == io_sinIndex[10:0] ? 30'h3e986a52 : _GEN_1221; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1223 = 11'hc6 == io_sinIndex[10:0] ? 30'h3e992a45 : _GEN_1222; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1224 = 11'hc7 == io_sinIndex[10:0] ? 30'h3e99ea1f : _GEN_1223; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1225 = 11'hc8 == io_sinIndex[10:0] ? 30'h3e9aa9e3 : _GEN_1224; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1226 = 11'hc9 == io_sinIndex[10:0] ? 30'h3e9b698e : _GEN_1225; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1227 = 11'hca == io_sinIndex[10:0] ? 30'h3e9c2921 : _GEN_1226; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1228 = 11'hcb == io_sinIndex[10:0] ? 30'h3e9ce89c : _GEN_1227; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1229 = 11'hcc == io_sinIndex[10:0] ? 30'h3e9da7ff : _GEN_1228; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1230 = 11'hcd == io_sinIndex[10:0] ? 30'h3e9e674a : _GEN_1229; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1231 = 11'hce == io_sinIndex[10:0] ? 30'h3e9f267c : _GEN_1230; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1232 = 11'hcf == io_sinIndex[10:0] ? 30'h3e9fe596 : _GEN_1231; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1233 = 11'hd0 == io_sinIndex[10:0] ? 30'h3ea0a497 : _GEN_1232; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1234 = 11'hd1 == io_sinIndex[10:0] ? 30'h3ea1637f : _GEN_1233; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1235 = 11'hd2 == io_sinIndex[10:0] ? 30'h3ea2224f : _GEN_1234; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1236 = 11'hd3 == io_sinIndex[10:0] ? 30'h3ea2e105 : _GEN_1235; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1237 = 11'hd4 == io_sinIndex[10:0] ? 30'h3ea39fa2 : _GEN_1236; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1238 = 11'hd5 == io_sinIndex[10:0] ? 30'h3ea45e26 : _GEN_1237; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1239 = 11'hd6 == io_sinIndex[10:0] ? 30'h3ea51c91 : _GEN_1238; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1240 = 11'hd7 == io_sinIndex[10:0] ? 30'h3ea5dae2 : _GEN_1239; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1241 = 11'hd8 == io_sinIndex[10:0] ? 30'h3ea69919 : _GEN_1240; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1242 = 11'hd9 == io_sinIndex[10:0] ? 30'h3ea75737 : _GEN_1241; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1243 = 11'hda == io_sinIndex[10:0] ? 30'h3ea8153b : _GEN_1242; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1244 = 11'hdb == io_sinIndex[10:0] ? 30'h3ea8d325 : _GEN_1243; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1245 = 11'hdc == io_sinIndex[10:0] ? 30'h3ea990f5 : _GEN_1244; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1246 = 11'hdd == io_sinIndex[10:0] ? 30'h3eaa4eab : _GEN_1245; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1247 = 11'hde == io_sinIndex[10:0] ? 30'h3eab0c47 : _GEN_1246; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1248 = 11'hdf == io_sinIndex[10:0] ? 30'h3eabc9c8 : _GEN_1247; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1249 = 11'he0 == io_sinIndex[10:0] ? 30'h3eac872f : _GEN_1248; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1250 = 11'he1 == io_sinIndex[10:0] ? 30'h3ead447b : _GEN_1249; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1251 = 11'he2 == io_sinIndex[10:0] ? 30'h3eae01ac : _GEN_1250; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1252 = 11'he3 == io_sinIndex[10:0] ? 30'h3eaebec3 : _GEN_1251; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1253 = 11'he4 == io_sinIndex[10:0] ? 30'h3eaf7bbe : _GEN_1252; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1254 = 11'he5 == io_sinIndex[10:0] ? 30'h3eb0389e : _GEN_1253; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1255 = 11'he6 == io_sinIndex[10:0] ? 30'h3eb0f564 : _GEN_1254; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1256 = 11'he7 == io_sinIndex[10:0] ? 30'h3eb1b20e : _GEN_1255; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1257 = 11'he8 == io_sinIndex[10:0] ? 30'h3eb26e9c : _GEN_1256; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1258 = 11'he9 == io_sinIndex[10:0] ? 30'h3eb32b0f : _GEN_1257; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1259 = 11'hea == io_sinIndex[10:0] ? 30'h3eb3e767 : _GEN_1258; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1260 = 11'heb == io_sinIndex[10:0] ? 30'h3eb4a3a2 : _GEN_1259; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1261 = 11'hec == io_sinIndex[10:0] ? 30'h3eb55fc2 : _GEN_1260; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1262 = 11'hed == io_sinIndex[10:0] ? 30'h3eb61bc6 : _GEN_1261; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1263 = 11'hee == io_sinIndex[10:0] ? 30'h3eb6d7ad : _GEN_1262; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1264 = 11'hef == io_sinIndex[10:0] ? 30'h3eb79379 : _GEN_1263; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1265 = 11'hf0 == io_sinIndex[10:0] ? 30'h3eb84f28 : _GEN_1264; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1266 = 11'hf1 == io_sinIndex[10:0] ? 30'h3eb90abb : _GEN_1265; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1267 = 11'hf2 == io_sinIndex[10:0] ? 30'h3eb9c631 : _GEN_1266; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1268 = 11'hf3 == io_sinIndex[10:0] ? 30'h3eba818a : _GEN_1267; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1269 = 11'hf4 == io_sinIndex[10:0] ? 30'h3ebb3cc7 : _GEN_1268; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1270 = 11'hf5 == io_sinIndex[10:0] ? 30'h3ebbf7e7 : _GEN_1269; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1271 = 11'hf6 == io_sinIndex[10:0] ? 30'h3ebcb2ea : _GEN_1270; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1272 = 11'hf7 == io_sinIndex[10:0] ? 30'h3ebd6dcf : _GEN_1271; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1273 = 11'hf8 == io_sinIndex[10:0] ? 30'h3ebe2898 : _GEN_1272; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1274 = 11'hf9 == io_sinIndex[10:0] ? 30'h3ebee343 : _GEN_1273; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1275 = 11'hfa == io_sinIndex[10:0] ? 30'h3ebf9dd1 : _GEN_1274; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1276 = 11'hfb == io_sinIndex[10:0] ? 30'h3ec05841 : _GEN_1275; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1277 = 11'hfc == io_sinIndex[10:0] ? 30'h3ec11293 : _GEN_1276; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1278 = 11'hfd == io_sinIndex[10:0] ? 30'h3ec1ccc8 : _GEN_1277; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1279 = 11'hfe == io_sinIndex[10:0] ? 30'h3ec286df : _GEN_1278; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1280 = 11'hff == io_sinIndex[10:0] ? 30'h3ec340d7 : _GEN_1279; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1281 = 11'h100 == io_sinIndex[10:0] ? 30'h3ec3fab2 : _GEN_1280; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1282 = 11'h101 == io_sinIndex[10:0] ? 30'h3ec4b46e : _GEN_1281; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1283 = 11'h102 == io_sinIndex[10:0] ? 30'h3ec56e0c : _GEN_1282; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1284 = 11'h103 == io_sinIndex[10:0] ? 30'h3ec6278c : _GEN_1283; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1285 = 11'h104 == io_sinIndex[10:0] ? 30'h3ec6e0ed : _GEN_1284; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1286 = 11'h105 == io_sinIndex[10:0] ? 30'h3ec79a2f : _GEN_1285; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1287 = 11'h106 == io_sinIndex[10:0] ? 30'h3ec85353 : _GEN_1286; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1288 = 11'h107 == io_sinIndex[10:0] ? 30'h3ec90c57 : _GEN_1287; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1289 = 11'h108 == io_sinIndex[10:0] ? 30'h3ec9c53d : _GEN_1288; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1290 = 11'h109 == io_sinIndex[10:0] ? 30'h3eca7e03 : _GEN_1289; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1291 = 11'h10a == io_sinIndex[10:0] ? 30'h3ecb36ab : _GEN_1290; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1292 = 11'h10b == io_sinIndex[10:0] ? 30'h3ecbef33 : _GEN_1291; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1293 = 11'h10c == io_sinIndex[10:0] ? 30'h3ecca79b : _GEN_1292; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1294 = 11'h10d == io_sinIndex[10:0] ? 30'h3ecd5fe4 : _GEN_1293; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1295 = 11'h10e == io_sinIndex[10:0] ? 30'h3ece180d : _GEN_1294; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1296 = 11'h10f == io_sinIndex[10:0] ? 30'h3eced016 : _GEN_1295; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1297 = 11'h110 == io_sinIndex[10:0] ? 30'h3ecf8800 : _GEN_1296; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1298 = 11'h111 == io_sinIndex[10:0] ? 30'h3ed03fc9 : _GEN_1297; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1299 = 11'h112 == io_sinIndex[10:0] ? 30'h3ed0f772 : _GEN_1298; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1300 = 11'h113 == io_sinIndex[10:0] ? 30'h3ed1aefb : _GEN_1299; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1301 = 11'h114 == io_sinIndex[10:0] ? 30'h3ed26664 : _GEN_1300; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1302 = 11'h115 == io_sinIndex[10:0] ? 30'h3ed31dac : _GEN_1301; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1303 = 11'h116 == io_sinIndex[10:0] ? 30'h3ed3d4d4 : _GEN_1302; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1304 = 11'h117 == io_sinIndex[10:0] ? 30'h3ed48bdb : _GEN_1303; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1305 = 11'h118 == io_sinIndex[10:0] ? 30'h3ed542c1 : _GEN_1304; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1306 = 11'h119 == io_sinIndex[10:0] ? 30'h3ed5f986 : _GEN_1305; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1307 = 11'h11a == io_sinIndex[10:0] ? 30'h3ed6b02b : _GEN_1306; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1308 = 11'h11b == io_sinIndex[10:0] ? 30'h3ed766ae : _GEN_1307; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1309 = 11'h11c == io_sinIndex[10:0] ? 30'h3ed81d10 : _GEN_1308; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1310 = 11'h11d == io_sinIndex[10:0] ? 30'h3ed8d350 : _GEN_1309; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1311 = 11'h11e == io_sinIndex[10:0] ? 30'h3ed9896f : _GEN_1310; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1312 = 11'h11f == io_sinIndex[10:0] ? 30'h3eda3f6d : _GEN_1311; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1313 = 11'h120 == io_sinIndex[10:0] ? 30'h3edaf549 : _GEN_1312; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1314 = 11'h121 == io_sinIndex[10:0] ? 30'h3edbab03 : _GEN_1313; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1315 = 11'h122 == io_sinIndex[10:0] ? 30'h3edc609b : _GEN_1314; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1316 = 11'h123 == io_sinIndex[10:0] ? 30'h3edd1611 : _GEN_1315; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1317 = 11'h124 == io_sinIndex[10:0] ? 30'h3eddcb65 : _GEN_1316; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1318 = 11'h125 == io_sinIndex[10:0] ? 30'h3ede8097 : _GEN_1317; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1319 = 11'h126 == io_sinIndex[10:0] ? 30'h3edf35a7 : _GEN_1318; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1320 = 11'h127 == io_sinIndex[10:0] ? 30'h3edfea94 : _GEN_1319; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1321 = 11'h128 == io_sinIndex[10:0] ? 30'h3ee09f5e : _GEN_1320; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1322 = 11'h129 == io_sinIndex[10:0] ? 30'h3ee15406 : _GEN_1321; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1323 = 11'h12a == io_sinIndex[10:0] ? 30'h3ee2088b : _GEN_1322; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1324 = 11'h12b == io_sinIndex[10:0] ? 30'h3ee2bced : _GEN_1323; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1325 = 11'h12c == io_sinIndex[10:0] ? 30'h3ee3712d : _GEN_1324; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1326 = 11'h12d == io_sinIndex[10:0] ? 30'h3ee42549 : _GEN_1325; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1327 = 11'h12e == io_sinIndex[10:0] ? 30'h3ee4d942 : _GEN_1326; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1328 = 11'h12f == io_sinIndex[10:0] ? 30'h3ee58d18 : _GEN_1327; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1329 = 11'h130 == io_sinIndex[10:0] ? 30'h3ee640ca : _GEN_1328; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1330 = 11'h131 == io_sinIndex[10:0] ? 30'h3ee6f459 : _GEN_1329; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1331 = 11'h132 == io_sinIndex[10:0] ? 30'h3ee7a7c4 : _GEN_1330; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1332 = 11'h133 == io_sinIndex[10:0] ? 30'h3ee85b0b : _GEN_1331; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1333 = 11'h134 == io_sinIndex[10:0] ? 30'h3ee90e2e : _GEN_1332; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1334 = 11'h135 == io_sinIndex[10:0] ? 30'h3ee9c12e : _GEN_1333; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1335 = 11'h136 == io_sinIndex[10:0] ? 30'h3eea7409 : _GEN_1334; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1336 = 11'h137 == io_sinIndex[10:0] ? 30'h3eeb26c1 : _GEN_1335; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1337 = 11'h138 == io_sinIndex[10:0] ? 30'h3eebd954 : _GEN_1336; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1338 = 11'h139 == io_sinIndex[10:0] ? 30'h3eec8bc2 : _GEN_1337; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1339 = 11'h13a == io_sinIndex[10:0] ? 30'h3eed3e0d : _GEN_1338; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1340 = 11'h13b == io_sinIndex[10:0] ? 30'h3eedf032 : _GEN_1339; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1341 = 11'h13c == io_sinIndex[10:0] ? 30'h3eeea233 : _GEN_1340; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1342 = 11'h13d == io_sinIndex[10:0] ? 30'h3eef540f : _GEN_1341; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1343 = 11'h13e == io_sinIndex[10:0] ? 30'h3ef005c6 : _GEN_1342; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1344 = 11'h13f == io_sinIndex[10:0] ? 30'h3ef0b758 : _GEN_1343; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1345 = 11'h140 == io_sinIndex[10:0] ? 30'h3ef168c5 : _GEN_1344; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1346 = 11'h141 == io_sinIndex[10:0] ? 30'h3ef21a0d : _GEN_1345; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1347 = 11'h142 == io_sinIndex[10:0] ? 30'h3ef2cb2f : _GEN_1346; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1348 = 11'h143 == io_sinIndex[10:0] ? 30'h3ef37c2c : _GEN_1347; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1349 = 11'h144 == io_sinIndex[10:0] ? 30'h3ef42d03 : _GEN_1348; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1350 = 11'h145 == io_sinIndex[10:0] ? 30'h3ef4ddb5 : _GEN_1349; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1351 = 11'h146 == io_sinIndex[10:0] ? 30'h3ef58e40 : _GEN_1350; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1352 = 11'h147 == io_sinIndex[10:0] ? 30'h3ef63ea6 : _GEN_1351; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1353 = 11'h148 == io_sinIndex[10:0] ? 30'h3ef6eee6 : _GEN_1352; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1354 = 11'h149 == io_sinIndex[10:0] ? 30'h3ef79f00 : _GEN_1353; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1355 = 11'h14a == io_sinIndex[10:0] ? 30'h3ef84ef4 : _GEN_1354; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1356 = 11'h14b == io_sinIndex[10:0] ? 30'h3ef8fec1 : _GEN_1355; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1357 = 11'h14c == io_sinIndex[10:0] ? 30'h3ef9ae68 : _GEN_1356; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1358 = 11'h14d == io_sinIndex[10:0] ? 30'h3efa5de8 : _GEN_1357; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1359 = 11'h14e == io_sinIndex[10:0] ? 30'h3efb0d42 : _GEN_1358; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1360 = 11'h14f == io_sinIndex[10:0] ? 30'h3efbbc75 : _GEN_1359; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1361 = 11'h150 == io_sinIndex[10:0] ? 30'h3efc6b81 : _GEN_1360; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1362 = 11'h151 == io_sinIndex[10:0] ? 30'h3efd1a67 : _GEN_1361; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1363 = 11'h152 == io_sinIndex[10:0] ? 30'h3efdc925 : _GEN_1362; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1364 = 11'h153 == io_sinIndex[10:0] ? 30'h3efe77bc : _GEN_1363; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1365 = 11'h154 == io_sinIndex[10:0] ? 30'h3eff262c : _GEN_1364; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1366 = 11'h155 == io_sinIndex[10:0] ? 30'h3effd474 : _GEN_1365; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1367 = 11'h156 == io_sinIndex[10:0] ? 30'h3f00414a : _GEN_1366; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1368 = 11'h157 == io_sinIndex[10:0] ? 30'h3f009847 : _GEN_1367; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1369 = 11'h158 == io_sinIndex[10:0] ? 30'h3f00ef30 : _GEN_1368; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1370 = 11'h159 == io_sinIndex[10:0] ? 30'h3f014605 : _GEN_1369; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1371 = 11'h15a == io_sinIndex[10:0] ? 30'h3f019cc6 : _GEN_1370; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1372 = 11'h15b == io_sinIndex[10:0] ? 30'h3f01f373 : _GEN_1371; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1373 = 11'h15c == io_sinIndex[10:0] ? 30'h3f024a0c : _GEN_1372; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1374 = 11'h15d == io_sinIndex[10:0] ? 30'h3f02a091 : _GEN_1373; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1375 = 11'h15e == io_sinIndex[10:0] ? 30'h3f02f701 : _GEN_1374; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1376 = 11'h15f == io_sinIndex[10:0] ? 30'h3f034d5e : _GEN_1375; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1377 = 11'h160 == io_sinIndex[10:0] ? 30'h3f03a3a6 : _GEN_1376; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1378 = 11'h161 == io_sinIndex[10:0] ? 30'h3f03f9da : _GEN_1377; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1379 = 11'h162 == io_sinIndex[10:0] ? 30'h3f044ffa : _GEN_1378; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1380 = 11'h163 == io_sinIndex[10:0] ? 30'h3f04a605 : _GEN_1379; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1381 = 11'h164 == io_sinIndex[10:0] ? 30'h3f04fbfc : _GEN_1380; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1382 = 11'h165 == io_sinIndex[10:0] ? 30'h3f0551de : _GEN_1381; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1383 = 11'h166 == io_sinIndex[10:0] ? 30'h3f05a7ab : _GEN_1382; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1384 = 11'h167 == io_sinIndex[10:0] ? 30'h3f05fd64 : _GEN_1383; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1385 = 11'h168 == io_sinIndex[10:0] ? 30'h3f065309 : _GEN_1384; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1386 = 11'h169 == io_sinIndex[10:0] ? 30'h3f06a898 : _GEN_1385; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1387 = 11'h16a == io_sinIndex[10:0] ? 30'h3f06fe13 : _GEN_1386; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1388 = 11'h16b == io_sinIndex[10:0] ? 30'h3f075379 : _GEN_1387; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1389 = 11'h16c == io_sinIndex[10:0] ? 30'h3f07a8ca : _GEN_1388; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1390 = 11'h16d == io_sinIndex[10:0] ? 30'h3f07fe06 : _GEN_1389; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1391 = 11'h16e == io_sinIndex[10:0] ? 30'h3f08532d : _GEN_1390; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1392 = 11'h16f == io_sinIndex[10:0] ? 30'h3f08a83f : _GEN_1391; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1393 = 11'h170 == io_sinIndex[10:0] ? 30'h3f08fd3d : _GEN_1392; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1394 = 11'h171 == io_sinIndex[10:0] ? 30'h3f095224 : _GEN_1393; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1395 = 11'h172 == io_sinIndex[10:0] ? 30'h3f09a6f7 : _GEN_1394; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1396 = 11'h173 == io_sinIndex[10:0] ? 30'h3f09fbb5 : _GEN_1395; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1397 = 11'h174 == io_sinIndex[10:0] ? 30'h3f0a505d : _GEN_1396; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1398 = 11'h175 == io_sinIndex[10:0] ? 30'h3f0aa4f0 : _GEN_1397; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1399 = 11'h176 == io_sinIndex[10:0] ? 30'h3f0af96d : _GEN_1398; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1400 = 11'h177 == io_sinIndex[10:0] ? 30'h3f0b4dd5 : _GEN_1399; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1401 = 11'h178 == io_sinIndex[10:0] ? 30'h3f0ba228 : _GEN_1400; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1402 = 11'h179 == io_sinIndex[10:0] ? 30'h3f0bf665 : _GEN_1401; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1403 = 11'h17a == io_sinIndex[10:0] ? 30'h3f0c4a8c : _GEN_1402; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1404 = 11'h17b == io_sinIndex[10:0] ? 30'h3f0c9e9e : _GEN_1403; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1405 = 11'h17c == io_sinIndex[10:0] ? 30'h3f0cf29a : _GEN_1404; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1406 = 11'h17d == io_sinIndex[10:0] ? 30'h3f0d4680 : _GEN_1405; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1407 = 11'h17e == io_sinIndex[10:0] ? 30'h3f0d9a51 : _GEN_1406; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1408 = 11'h17f == io_sinIndex[10:0] ? 30'h3f0dee0c : _GEN_1407; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1409 = 11'h180 == io_sinIndex[10:0] ? 30'h3f0e41b0 : _GEN_1408; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1410 = 11'h181 == io_sinIndex[10:0] ? 30'h3f0e953f : _GEN_1409; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1411 = 11'h182 == io_sinIndex[10:0] ? 30'h3f0ee8b8 : _GEN_1410; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1412 = 11'h183 == io_sinIndex[10:0] ? 30'h3f0f3c1b : _GEN_1411; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1413 = 11'h184 == io_sinIndex[10:0] ? 30'h3f0f8f67 : _GEN_1412; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1414 = 11'h185 == io_sinIndex[10:0] ? 30'h3f0fe29e : _GEN_1413; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1415 = 11'h186 == io_sinIndex[10:0] ? 30'h3f1035be : _GEN_1414; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1416 = 11'h187 == io_sinIndex[10:0] ? 30'h3f1088c8 : _GEN_1415; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1417 = 11'h188 == io_sinIndex[10:0] ? 30'h3f10dbbc : _GEN_1416; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1418 = 11'h189 == io_sinIndex[10:0] ? 30'h3f112e9a : _GEN_1417; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1419 = 11'h18a == io_sinIndex[10:0] ? 30'h3f118161 : _GEN_1418; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1420 = 11'h18b == io_sinIndex[10:0] ? 30'h3f11d411 : _GEN_1419; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1421 = 11'h18c == io_sinIndex[10:0] ? 30'h3f1226ab : _GEN_1420; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1422 = 11'h18d == io_sinIndex[10:0] ? 30'h3f12792f : _GEN_1421; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1423 = 11'h18e == io_sinIndex[10:0] ? 30'h3f12cb9c : _GEN_1422; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1424 = 11'h18f == io_sinIndex[10:0] ? 30'h3f131df2 : _GEN_1423; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1425 = 11'h190 == io_sinIndex[10:0] ? 30'h3f137032 : _GEN_1424; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1426 = 11'h191 == io_sinIndex[10:0] ? 30'h3f13c25a : _GEN_1425; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1427 = 11'h192 == io_sinIndex[10:0] ? 30'h3f14146c : _GEN_1426; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1428 = 11'h193 == io_sinIndex[10:0] ? 30'h3f146668 : _GEN_1427; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1429 = 11'h194 == io_sinIndex[10:0] ? 30'h3f14b84c : _GEN_1428; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1430 = 11'h195 == io_sinIndex[10:0] ? 30'h3f150a19 : _GEN_1429; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1431 = 11'h196 == io_sinIndex[10:0] ? 30'h3f155bd0 : _GEN_1430; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1432 = 11'h197 == io_sinIndex[10:0] ? 30'h3f15ad6f : _GEN_1431; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1433 = 11'h198 == io_sinIndex[10:0] ? 30'h3f15fef7 : _GEN_1432; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1434 = 11'h199 == io_sinIndex[10:0] ? 30'h3f165068 : _GEN_1433; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1435 = 11'h19a == io_sinIndex[10:0] ? 30'h3f16a1c2 : _GEN_1434; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1436 = 11'h19b == io_sinIndex[10:0] ? 30'h3f16f305 : _GEN_1435; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1437 = 11'h19c == io_sinIndex[10:0] ? 30'h3f174430 : _GEN_1436; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1438 = 11'h19d == io_sinIndex[10:0] ? 30'h3f179544 : _GEN_1437; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1439 = 11'h19e == io_sinIndex[10:0] ? 30'h3f17e641 : _GEN_1438; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1440 = 11'h19f == io_sinIndex[10:0] ? 30'h3f183726 : _GEN_1439; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1441 = 11'h1a0 == io_sinIndex[10:0] ? 30'h3f1887f4 : _GEN_1440; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1442 = 11'h1a1 == io_sinIndex[10:0] ? 30'h3f18d8aa : _GEN_1441; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1443 = 11'h1a2 == io_sinIndex[10:0] ? 30'h3f192948 : _GEN_1442; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1444 = 11'h1a3 == io_sinIndex[10:0] ? 30'h3f1979cf : _GEN_1443; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1445 = 11'h1a4 == io_sinIndex[10:0] ? 30'h3f19ca3f : _GEN_1444; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1446 = 11'h1a5 == io_sinIndex[10:0] ? 30'h3f1a1a96 : _GEN_1445; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1447 = 11'h1a6 == io_sinIndex[10:0] ? 30'h3f1a6ad6 : _GEN_1446; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1448 = 11'h1a7 == io_sinIndex[10:0] ? 30'h3f1abafe : _GEN_1447; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1449 = 11'h1a8 == io_sinIndex[10:0] ? 30'h3f1b0b0e : _GEN_1448; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1450 = 11'h1a9 == io_sinIndex[10:0] ? 30'h3f1b5b06 : _GEN_1449; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1451 = 11'h1aa == io_sinIndex[10:0] ? 30'h3f1baae6 : _GEN_1450; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1452 = 11'h1ab == io_sinIndex[10:0] ? 30'h3f1bfaaf : _GEN_1451; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1453 = 11'h1ac == io_sinIndex[10:0] ? 30'h3f1c4a5f : _GEN_1452; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1454 = 11'h1ad == io_sinIndex[10:0] ? 30'h3f1c99f7 : _GEN_1453; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1455 = 11'h1ae == io_sinIndex[10:0] ? 30'h3f1ce977 : _GEN_1454; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1456 = 11'h1af == io_sinIndex[10:0] ? 30'h3f1d38de : _GEN_1455; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1457 = 11'h1b0 == io_sinIndex[10:0] ? 30'h3f1d882e : _GEN_1456; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1458 = 11'h1b1 == io_sinIndex[10:0] ? 30'h3f1dd765 : _GEN_1457; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1459 = 11'h1b2 == io_sinIndex[10:0] ? 30'h3f1e2683 : _GEN_1458; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1460 = 11'h1b3 == io_sinIndex[10:0] ? 30'h3f1e758a : _GEN_1459; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1461 = 11'h1b4 == io_sinIndex[10:0] ? 30'h3f1ec477 : _GEN_1460; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1462 = 11'h1b5 == io_sinIndex[10:0] ? 30'h3f1f134d : _GEN_1461; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1463 = 11'h1b6 == io_sinIndex[10:0] ? 30'h3f1f620a : _GEN_1462; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1464 = 11'h1b7 == io_sinIndex[10:0] ? 30'h3f1fb0ae : _GEN_1463; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1465 = 11'h1b8 == io_sinIndex[10:0] ? 30'h3f1fff39 : _GEN_1464; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1466 = 11'h1b9 == io_sinIndex[10:0] ? 30'h3f204dac : _GEN_1465; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1467 = 11'h1ba == io_sinIndex[10:0] ? 30'h3f209c06 : _GEN_1466; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1468 = 11'h1bb == io_sinIndex[10:0] ? 30'h3f20ea48 : _GEN_1467; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1469 = 11'h1bc == io_sinIndex[10:0] ? 30'h3f213870 : _GEN_1468; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1470 = 11'h1bd == io_sinIndex[10:0] ? 30'h3f218680 : _GEN_1469; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1471 = 11'h1be == io_sinIndex[10:0] ? 30'h3f21d477 : _GEN_1470; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1472 = 11'h1bf == io_sinIndex[10:0] ? 30'h3f222255 : _GEN_1471; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1473 = 11'h1c0 == io_sinIndex[10:0] ? 30'h3f227019 : _GEN_1472; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1474 = 11'h1c1 == io_sinIndex[10:0] ? 30'h3f22bdc5 : _GEN_1473; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1475 = 11'h1c2 == io_sinIndex[10:0] ? 30'h3f230b58 : _GEN_1474; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1476 = 11'h1c3 == io_sinIndex[10:0] ? 30'h3f2358d1 : _GEN_1475; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1477 = 11'h1c4 == io_sinIndex[10:0] ? 30'h3f23a631 : _GEN_1476; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1478 = 11'h1c5 == io_sinIndex[10:0] ? 30'h3f23f378 : _GEN_1477; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1479 = 11'h1c6 == io_sinIndex[10:0] ? 30'h3f2440a6 : _GEN_1478; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1480 = 11'h1c7 == io_sinIndex[10:0] ? 30'h3f248dbb : _GEN_1479; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1481 = 11'h1c8 == io_sinIndex[10:0] ? 30'h3f24dab6 : _GEN_1480; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1482 = 11'h1c9 == io_sinIndex[10:0] ? 30'h3f252797 : _GEN_1481; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1483 = 11'h1ca == io_sinIndex[10:0] ? 30'h3f25745f : _GEN_1482; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1484 = 11'h1cb == io_sinIndex[10:0] ? 30'h3f25c10e : _GEN_1483; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1485 = 11'h1cc == io_sinIndex[10:0] ? 30'h3f260da3 : _GEN_1484; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1486 = 11'h1cd == io_sinIndex[10:0] ? 30'h3f265a1e : _GEN_1485; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1487 = 11'h1ce == io_sinIndex[10:0] ? 30'h3f26a680 : _GEN_1486; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1488 = 11'h1cf == io_sinIndex[10:0] ? 30'h3f26f2c8 : _GEN_1487; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1489 = 11'h1d0 == io_sinIndex[10:0] ? 30'h3f273ef6 : _GEN_1488; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1490 = 11'h1d1 == io_sinIndex[10:0] ? 30'h3f278b0a : _GEN_1489; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1491 = 11'h1d2 == io_sinIndex[10:0] ? 30'h3f27d705 : _GEN_1490; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1492 = 11'h1d3 == io_sinIndex[10:0] ? 30'h3f2822e5 : _GEN_1491; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1493 = 11'h1d4 == io_sinIndex[10:0] ? 30'h3f286eac : _GEN_1492; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1494 = 11'h1d5 == io_sinIndex[10:0] ? 30'h3f28ba59 : _GEN_1493; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1495 = 11'h1d6 == io_sinIndex[10:0] ? 30'h3f2905ec : _GEN_1494; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1496 = 11'h1d7 == io_sinIndex[10:0] ? 30'h3f295164 : _GEN_1495; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1497 = 11'h1d8 == io_sinIndex[10:0] ? 30'h3f299cc3 : _GEN_1496; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1498 = 11'h1d9 == io_sinIndex[10:0] ? 30'h3f29e807 : _GEN_1497; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1499 = 11'h1da == io_sinIndex[10:0] ? 30'h3f2a3331 : _GEN_1498; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1500 = 11'h1db == io_sinIndex[10:0] ? 30'h3f2a7e41 : _GEN_1499; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1501 = 11'h1dc == io_sinIndex[10:0] ? 30'h3f2ac936 : _GEN_1500; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1502 = 11'h1dd == io_sinIndex[10:0] ? 30'h3f2b1412 : _GEN_1501; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1503 = 11'h1de == io_sinIndex[10:0] ? 30'h3f2b5ed2 : _GEN_1502; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1504 = 11'h1df == io_sinIndex[10:0] ? 30'h3f2ba979 : _GEN_1503; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1505 = 11'h1e0 == io_sinIndex[10:0] ? 30'h3f2bf405 : _GEN_1504; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1506 = 11'h1e1 == io_sinIndex[10:0] ? 30'h3f2c3e76 : _GEN_1505; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1507 = 11'h1e2 == io_sinIndex[10:0] ? 30'h3f2c88cd : _GEN_1506; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1508 = 11'h1e3 == io_sinIndex[10:0] ? 30'h3f2cd309 : _GEN_1507; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1509 = 11'h1e4 == io_sinIndex[10:0] ? 30'h3f2d1d2a : _GEN_1508; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1510 = 11'h1e5 == io_sinIndex[10:0] ? 30'h3f2d6731 : _GEN_1509; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1511 = 11'h1e6 == io_sinIndex[10:0] ? 30'h3f2db11d : _GEN_1510; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1512 = 11'h1e7 == io_sinIndex[10:0] ? 30'h3f2dfaee : _GEN_1511; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1513 = 11'h1e8 == io_sinIndex[10:0] ? 30'h3f2e44a5 : _GEN_1512; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1514 = 11'h1e9 == io_sinIndex[10:0] ? 30'h3f2e8e40 : _GEN_1513; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1515 = 11'h1ea == io_sinIndex[10:0] ? 30'h3f2ed7c1 : _GEN_1514; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1516 = 11'h1eb == io_sinIndex[10:0] ? 30'h3f2f2126 : _GEN_1515; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1517 = 11'h1ec == io_sinIndex[10:0] ? 30'h3f2f6a71 : _GEN_1516; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1518 = 11'h1ed == io_sinIndex[10:0] ? 30'h3f2fb3a0 : _GEN_1517; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1519 = 11'h1ee == io_sinIndex[10:0] ? 30'h3f2ffcb5 : _GEN_1518; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1520 = 11'h1ef == io_sinIndex[10:0] ? 30'h3f3045ae : _GEN_1519; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1521 = 11'h1f0 == io_sinIndex[10:0] ? 30'h3f308e8c : _GEN_1520; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1522 = 11'h1f1 == io_sinIndex[10:0] ? 30'h3f30d74f : _GEN_1521; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1523 = 11'h1f2 == io_sinIndex[10:0] ? 30'h3f311ff6 : _GEN_1522; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1524 = 11'h1f3 == io_sinIndex[10:0] ? 30'h3f316883 : _GEN_1523; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1525 = 11'h1f4 == io_sinIndex[10:0] ? 30'h3f31b0f3 : _GEN_1524; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1526 = 11'h1f5 == io_sinIndex[10:0] ? 30'h3f31f949 : _GEN_1525; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1527 = 11'h1f6 == io_sinIndex[10:0] ? 30'h3f324183 : _GEN_1526; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1528 = 11'h1f7 == io_sinIndex[10:0] ? 30'h3f3289a1 : _GEN_1527; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1529 = 11'h1f8 == io_sinIndex[10:0] ? 30'h3f32d1a4 : _GEN_1528; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1530 = 11'h1f9 == io_sinIndex[10:0] ? 30'h3f33198b : _GEN_1529; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1531 = 11'h1fa == io_sinIndex[10:0] ? 30'h3f336157 : _GEN_1530; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1532 = 11'h1fb == io_sinIndex[10:0] ? 30'h3f33a907 : _GEN_1531; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1533 = 11'h1fc == io_sinIndex[10:0] ? 30'h3f33f09b : _GEN_1532; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1534 = 11'h1fd == io_sinIndex[10:0] ? 30'h3f343814 : _GEN_1533; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1535 = 11'h1fe == io_sinIndex[10:0] ? 30'h3f347f70 : _GEN_1534; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1536 = 11'h1ff == io_sinIndex[10:0] ? 30'h3f34c6b1 : _GEN_1535; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1537 = 11'h200 == io_sinIndex[10:0] ? 30'h3f350dd6 : _GEN_1536; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1538 = 11'h201 == io_sinIndex[10:0] ? 30'h3f3554df : _GEN_1537; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1539 = 11'h202 == io_sinIndex[10:0] ? 30'h3f359bcc : _GEN_1538; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1540 = 11'h203 == io_sinIndex[10:0] ? 30'h3f35e29d : _GEN_1539; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1541 = 11'h204 == io_sinIndex[10:0] ? 30'h3f362952 : _GEN_1540; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1542 = 11'h205 == io_sinIndex[10:0] ? 30'h3f366feb : _GEN_1541; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1543 = 11'h206 == io_sinIndex[10:0] ? 30'h3f36b668 : _GEN_1542; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1544 = 11'h207 == io_sinIndex[10:0] ? 30'h3f36fcc8 : _GEN_1543; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1545 = 11'h208 == io_sinIndex[10:0] ? 30'h3f37430d : _GEN_1544; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1546 = 11'h209 == io_sinIndex[10:0] ? 30'h3f378935 : _GEN_1545; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1547 = 11'h20a == io_sinIndex[10:0] ? 30'h3f37cf40 : _GEN_1546; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1548 = 11'h20b == io_sinIndex[10:0] ? 30'h3f381530 : _GEN_1547; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1549 = 11'h20c == io_sinIndex[10:0] ? 30'h3f385b03 : _GEN_1548; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1550 = 11'h20d == io_sinIndex[10:0] ? 30'h3f38a0b9 : _GEN_1549; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1551 = 11'h20e == io_sinIndex[10:0] ? 30'h3f38e653 : _GEN_1550; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1552 = 11'h20f == io_sinIndex[10:0] ? 30'h3f392bd1 : _GEN_1551; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1553 = 11'h210 == io_sinIndex[10:0] ? 30'h3f397132 : _GEN_1552; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1554 = 11'h211 == io_sinIndex[10:0] ? 30'h3f39b676 : _GEN_1553; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1555 = 11'h212 == io_sinIndex[10:0] ? 30'h3f39fb9e : _GEN_1554; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1556 = 11'h213 == io_sinIndex[10:0] ? 30'h3f3a40a9 : _GEN_1555; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1557 = 11'h214 == io_sinIndex[10:0] ? 30'h3f3a8597 : _GEN_1556; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1558 = 11'h215 == io_sinIndex[10:0] ? 30'h3f3aca68 : _GEN_1557; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1559 = 11'h216 == io_sinIndex[10:0] ? 30'h3f3b0f1d : _GEN_1558; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1560 = 11'h217 == io_sinIndex[10:0] ? 30'h3f3b53b5 : _GEN_1559; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1561 = 11'h218 == io_sinIndex[10:0] ? 30'h3f3b982f : _GEN_1560; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1562 = 11'h219 == io_sinIndex[10:0] ? 30'h3f3bdc8d : _GEN_1561; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1563 = 11'h21a == io_sinIndex[10:0] ? 30'h3f3c20ce : _GEN_1562; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1564 = 11'h21b == io_sinIndex[10:0] ? 30'h3f3c64f2 : _GEN_1563; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1565 = 11'h21c == io_sinIndex[10:0] ? 30'h3f3ca8f9 : _GEN_1564; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1566 = 11'h21d == io_sinIndex[10:0] ? 30'h3f3cece3 : _GEN_1565; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1567 = 11'h21e == io_sinIndex[10:0] ? 30'h3f3d30af : _GEN_1566; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1568 = 11'h21f == io_sinIndex[10:0] ? 30'h3f3d745f : _GEN_1567; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1569 = 11'h220 == io_sinIndex[10:0] ? 30'h3f3db7f1 : _GEN_1568; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1570 = 11'h221 == io_sinIndex[10:0] ? 30'h3f3dfb66 : _GEN_1569; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1571 = 11'h222 == io_sinIndex[10:0] ? 30'h3f3e3ebd : _GEN_1570; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1572 = 11'h223 == io_sinIndex[10:0] ? 30'h3f3e81f7 : _GEN_1571; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1573 = 11'h224 == io_sinIndex[10:0] ? 30'h3f3ec514 : _GEN_1572; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1574 = 11'h225 == io_sinIndex[10:0] ? 30'h3f3f0814 : _GEN_1573; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1575 = 11'h226 == io_sinIndex[10:0] ? 30'h3f3f4af6 : _GEN_1574; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1576 = 11'h227 == io_sinIndex[10:0] ? 30'h3f3f8dba : _GEN_1575; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1577 = 11'h228 == io_sinIndex[10:0] ? 30'h3f3fd061 : _GEN_1576; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1578 = 11'h229 == io_sinIndex[10:0] ? 30'h3f4012ea : _GEN_1577; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1579 = 11'h22a == io_sinIndex[10:0] ? 30'h3f405556 : _GEN_1578; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1580 = 11'h22b == io_sinIndex[10:0] ? 30'h3f4097a4 : _GEN_1579; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1581 = 11'h22c == io_sinIndex[10:0] ? 30'h3f40d9d4 : _GEN_1580; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1582 = 11'h22d == io_sinIndex[10:0] ? 30'h3f411be6 : _GEN_1581; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1583 = 11'h22e == io_sinIndex[10:0] ? 30'h3f415ddb : _GEN_1582; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1584 = 11'h22f == io_sinIndex[10:0] ? 30'h3f419fb2 : _GEN_1583; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1585 = 11'h230 == io_sinIndex[10:0] ? 30'h3f41e16b : _GEN_1584; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1586 = 11'h231 == io_sinIndex[10:0] ? 30'h3f422306 : _GEN_1585; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1587 = 11'h232 == io_sinIndex[10:0] ? 30'h3f426483 : _GEN_1586; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1588 = 11'h233 == io_sinIndex[10:0] ? 30'h3f42a5e2 : _GEN_1587; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1589 = 11'h234 == io_sinIndex[10:0] ? 30'h3f42e723 : _GEN_1588; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1590 = 11'h235 == io_sinIndex[10:0] ? 30'h3f432846 : _GEN_1589; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1591 = 11'h236 == io_sinIndex[10:0] ? 30'h3f43694b : _GEN_1590; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1592 = 11'h237 == io_sinIndex[10:0] ? 30'h3f43aa32 : _GEN_1591; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1593 = 11'h238 == io_sinIndex[10:0] ? 30'h3f43eafa : _GEN_1592; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1594 = 11'h239 == io_sinIndex[10:0] ? 30'h3f442ba5 : _GEN_1593; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1595 = 11'h23a == io_sinIndex[10:0] ? 30'h3f446c31 : _GEN_1594; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1596 = 11'h23b == io_sinIndex[10:0] ? 30'h3f44ac9f : _GEN_1595; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1597 = 11'h23c == io_sinIndex[10:0] ? 30'h3f44ecee : _GEN_1596; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1598 = 11'h23d == io_sinIndex[10:0] ? 30'h3f452d1f : _GEN_1597; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1599 = 11'h23e == io_sinIndex[10:0] ? 30'h3f456d32 : _GEN_1598; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1600 = 11'h23f == io_sinIndex[10:0] ? 30'h3f45ad26 : _GEN_1599; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1601 = 11'h240 == io_sinIndex[10:0] ? 30'h3f45ecfc : _GEN_1600; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1602 = 11'h241 == io_sinIndex[10:0] ? 30'h3f462cb3 : _GEN_1601; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1603 = 11'h242 == io_sinIndex[10:0] ? 30'h3f466c4b : _GEN_1602; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1604 = 11'h243 == io_sinIndex[10:0] ? 30'h3f46abc5 : _GEN_1603; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1605 = 11'h244 == io_sinIndex[10:0] ? 30'h3f46eb20 : _GEN_1604; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1606 = 11'h245 == io_sinIndex[10:0] ? 30'h3f472a5d : _GEN_1605; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1607 = 11'h246 == io_sinIndex[10:0] ? 30'h3f47697b : _GEN_1606; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1608 = 11'h247 == io_sinIndex[10:0] ? 30'h3f47a87a : _GEN_1607; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1609 = 11'h248 == io_sinIndex[10:0] ? 30'h3f47e75a : _GEN_1608; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1610 = 11'h249 == io_sinIndex[10:0] ? 30'h3f48261c : _GEN_1609; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1611 = 11'h24a == io_sinIndex[10:0] ? 30'h3f4864be : _GEN_1610; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1612 = 11'h24b == io_sinIndex[10:0] ? 30'h3f48a342 : _GEN_1611; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1613 = 11'h24c == io_sinIndex[10:0] ? 30'h3f48e1a7 : _GEN_1612; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1614 = 11'h24d == io_sinIndex[10:0] ? 30'h3f491fec : _GEN_1613; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1615 = 11'h24e == io_sinIndex[10:0] ? 30'h3f495e13 : _GEN_1614; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1616 = 11'h24f == io_sinIndex[10:0] ? 30'h3f499c1a : _GEN_1615; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1617 = 11'h250 == io_sinIndex[10:0] ? 30'h3f49da03 : _GEN_1616; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1618 = 11'h251 == io_sinIndex[10:0] ? 30'h3f4a17cc : _GEN_1617; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1619 = 11'h252 == io_sinIndex[10:0] ? 30'h3f4a5576 : _GEN_1618; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1620 = 11'h253 == io_sinIndex[10:0] ? 30'h3f4a9301 : _GEN_1619; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1621 = 11'h254 == io_sinIndex[10:0] ? 30'h3f4ad06d : _GEN_1620; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1622 = 11'h255 == io_sinIndex[10:0] ? 30'h3f4b0dba : _GEN_1621; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1623 = 11'h256 == io_sinIndex[10:0] ? 30'h3f4b4ae7 : _GEN_1622; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1624 = 11'h257 == io_sinIndex[10:0] ? 30'h3f4b87f4 : _GEN_1623; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1625 = 11'h258 == io_sinIndex[10:0] ? 30'h3f4bc4e3 : _GEN_1624; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1626 = 11'h259 == io_sinIndex[10:0] ? 30'h3f4c01b1 : _GEN_1625; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1627 = 11'h25a == io_sinIndex[10:0] ? 30'h3f4c3e61 : _GEN_1626; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1628 = 11'h25b == io_sinIndex[10:0] ? 30'h3f4c7af1 : _GEN_1627; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1629 = 11'h25c == io_sinIndex[10:0] ? 30'h3f4cb761 : _GEN_1628; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1630 = 11'h25d == io_sinIndex[10:0] ? 30'h3f4cf3b2 : _GEN_1629; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1631 = 11'h25e == io_sinIndex[10:0] ? 30'h3f4d2fe3 : _GEN_1630; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1632 = 11'h25f == io_sinIndex[10:0] ? 30'h3f4d6bf4 : _GEN_1631; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1633 = 11'h260 == io_sinIndex[10:0] ? 30'h3f4da7e6 : _GEN_1632; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1634 = 11'h261 == io_sinIndex[10:0] ? 30'h3f4de3b8 : _GEN_1633; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1635 = 11'h262 == io_sinIndex[10:0] ? 30'h3f4e1f6a : _GEN_1634; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1636 = 11'h263 == io_sinIndex[10:0] ? 30'h3f4e5afd : _GEN_1635; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1637 = 11'h264 == io_sinIndex[10:0] ? 30'h3f4e9670 : _GEN_1636; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1638 = 11'h265 == io_sinIndex[10:0] ? 30'h3f4ed1c2 : _GEN_1637; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1639 = 11'h266 == io_sinIndex[10:0] ? 30'h3f4f0cf5 : _GEN_1638; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1640 = 11'h267 == io_sinIndex[10:0] ? 30'h3f4f4808 : _GEN_1639; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1641 = 11'h268 == io_sinIndex[10:0] ? 30'h3f4f82fb : _GEN_1640; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1642 = 11'h269 == io_sinIndex[10:0] ? 30'h3f4fbdce : _GEN_1641; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1643 = 11'h26a == io_sinIndex[10:0] ? 30'h3f4ff881 : _GEN_1642; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1644 = 11'h26b == io_sinIndex[10:0] ? 30'h3f503313 : _GEN_1643; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1645 = 11'h26c == io_sinIndex[10:0] ? 30'h3f506d86 : _GEN_1644; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1646 = 11'h26d == io_sinIndex[10:0] ? 30'h3f50a7d9 : _GEN_1645; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1647 = 11'h26e == io_sinIndex[10:0] ? 30'h3f50e20b : _GEN_1646; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1648 = 11'h26f == io_sinIndex[10:0] ? 30'h3f511c1d : _GEN_1647; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1649 = 11'h270 == io_sinIndex[10:0] ? 30'h3f51560f : _GEN_1648; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1650 = 11'h271 == io_sinIndex[10:0] ? 30'h3f518fe0 : _GEN_1649; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1651 = 11'h272 == io_sinIndex[10:0] ? 30'h3f51c991 : _GEN_1650; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1652 = 11'h273 == io_sinIndex[10:0] ? 30'h3f520322 : _GEN_1651; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1653 = 11'h274 == io_sinIndex[10:0] ? 30'h3f523c93 : _GEN_1652; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1654 = 11'h275 == io_sinIndex[10:0] ? 30'h3f5275e3 : _GEN_1653; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1655 = 11'h276 == io_sinIndex[10:0] ? 30'h3f52af12 : _GEN_1654; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1656 = 11'h277 == io_sinIndex[10:0] ? 30'h3f52e821 : _GEN_1655; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1657 = 11'h278 == io_sinIndex[10:0] ? 30'h3f532110 : _GEN_1656; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1658 = 11'h279 == io_sinIndex[10:0] ? 30'h3f5359dd : _GEN_1657; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1659 = 11'h27a == io_sinIndex[10:0] ? 30'h3f53928b : _GEN_1658; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1660 = 11'h27b == io_sinIndex[10:0] ? 30'h3f53cb17 : _GEN_1659; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1661 = 11'h27c == io_sinIndex[10:0] ? 30'h3f540383 : _GEN_1660; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1662 = 11'h27d == io_sinIndex[10:0] ? 30'h3f543bce : _GEN_1661; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1663 = 11'h27e == io_sinIndex[10:0] ? 30'h3f5473f9 : _GEN_1662; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1664 = 11'h27f == io_sinIndex[10:0] ? 30'h3f54ac03 : _GEN_1663; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1665 = 11'h280 == io_sinIndex[10:0] ? 30'h3f54e3ec : _GEN_1664; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1666 = 11'h281 == io_sinIndex[10:0] ? 30'h3f551bb4 : _GEN_1665; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1667 = 11'h282 == io_sinIndex[10:0] ? 30'h3f55535b : _GEN_1666; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1668 = 11'h283 == io_sinIndex[10:0] ? 30'h3f558ae1 : _GEN_1667; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1669 = 11'h284 == io_sinIndex[10:0] ? 30'h3f55c246 : _GEN_1668; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1670 = 11'h285 == io_sinIndex[10:0] ? 30'h3f55f98b : _GEN_1669; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1671 = 11'h286 == io_sinIndex[10:0] ? 30'h3f5630ae : _GEN_1670; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1672 = 11'h287 == io_sinIndex[10:0] ? 30'h3f5667b0 : _GEN_1671; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1673 = 11'h288 == io_sinIndex[10:0] ? 30'h3f569e91 : _GEN_1672; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1674 = 11'h289 == io_sinIndex[10:0] ? 30'h3f56d551 : _GEN_1673; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1675 = 11'h28a == io_sinIndex[10:0] ? 30'h3f570bf0 : _GEN_1674; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1676 = 11'h28b == io_sinIndex[10:0] ? 30'h3f57426e : _GEN_1675; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1677 = 11'h28c == io_sinIndex[10:0] ? 30'h3f5778cb : _GEN_1676; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1678 = 11'h28d == io_sinIndex[10:0] ? 30'h3f57af06 : _GEN_1677; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1679 = 11'h28e == io_sinIndex[10:0] ? 30'h3f57e520 : _GEN_1678; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1680 = 11'h28f == io_sinIndex[10:0] ? 30'h3f581b19 : _GEN_1679; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1681 = 11'h290 == io_sinIndex[10:0] ? 30'h3f5850f0 : _GEN_1680; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1682 = 11'h291 == io_sinIndex[10:0] ? 30'h3f5886a6 : _GEN_1681; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1683 = 11'h292 == io_sinIndex[10:0] ? 30'h3f58bc3b : _GEN_1682; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1684 = 11'h293 == io_sinIndex[10:0] ? 30'h3f58f1ae : _GEN_1683; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1685 = 11'h294 == io_sinIndex[10:0] ? 30'h3f5926ff : _GEN_1684; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1686 = 11'h295 == io_sinIndex[10:0] ? 30'h3f595c30 : _GEN_1685; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1687 = 11'h296 == io_sinIndex[10:0] ? 30'h3f59913e : _GEN_1686; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1688 = 11'h297 == io_sinIndex[10:0] ? 30'h3f59c62b : _GEN_1687; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1689 = 11'h298 == io_sinIndex[10:0] ? 30'h3f59faf7 : _GEN_1688; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1690 = 11'h299 == io_sinIndex[10:0] ? 30'h3f5a2fa0 : _GEN_1689; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1691 = 11'h29a == io_sinIndex[10:0] ? 30'h3f5a6429 : _GEN_1690; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1692 = 11'h29b == io_sinIndex[10:0] ? 30'h3f5a988f : _GEN_1691; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1693 = 11'h29c == io_sinIndex[10:0] ? 30'h3f5accd4 : _GEN_1692; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1694 = 11'h29d == io_sinIndex[10:0] ? 30'h3f5b00f7 : _GEN_1693; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1695 = 11'h29e == io_sinIndex[10:0] ? 30'h3f5b34f8 : _GEN_1694; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1696 = 11'h29f == io_sinIndex[10:0] ? 30'h3f5b68d7 : _GEN_1695; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1697 = 11'h2a0 == io_sinIndex[10:0] ? 30'h3f5b9c95 : _GEN_1696; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1698 = 11'h2a1 == io_sinIndex[10:0] ? 30'h3f5bd031 : _GEN_1697; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1699 = 11'h2a2 == io_sinIndex[10:0] ? 30'h3f5c03aa : _GEN_1698; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1700 = 11'h2a3 == io_sinIndex[10:0] ? 30'h3f5c3702 : _GEN_1699; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1701 = 11'h2a4 == io_sinIndex[10:0] ? 30'h3f5c6a38 : _GEN_1700; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1702 = 11'h2a5 == io_sinIndex[10:0] ? 30'h3f5c9d4c : _GEN_1701; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1703 = 11'h2a6 == io_sinIndex[10:0] ? 30'h3f5cd03d : _GEN_1702; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1704 = 11'h2a7 == io_sinIndex[10:0] ? 30'h3f5d030d : _GEN_1703; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1705 = 11'h2a8 == io_sinIndex[10:0] ? 30'h3f5d35bb : _GEN_1704; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1706 = 11'h2a9 == io_sinIndex[10:0] ? 30'h3f5d6846 : _GEN_1705; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1707 = 11'h2aa == io_sinIndex[10:0] ? 30'h3f5d9aaf : _GEN_1706; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1708 = 11'h2ab == io_sinIndex[10:0] ? 30'h3f5dccf7 : _GEN_1707; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1709 = 11'h2ac == io_sinIndex[10:0] ? 30'h3f5dff1b : _GEN_1708; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1710 = 11'h2ad == io_sinIndex[10:0] ? 30'h3f5e311e : _GEN_1709; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1711 = 11'h2ae == io_sinIndex[10:0] ? 30'h3f5e62fe : _GEN_1710; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1712 = 11'h2af == io_sinIndex[10:0] ? 30'h3f5e94bc : _GEN_1711; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1713 = 11'h2b0 == io_sinIndex[10:0] ? 30'h3f5ec658 : _GEN_1712; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1714 = 11'h2b1 == io_sinIndex[10:0] ? 30'h3f5ef7d1 : _GEN_1713; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1715 = 11'h2b2 == io_sinIndex[10:0] ? 30'h3f5f2928 : _GEN_1714; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1716 = 11'h2b3 == io_sinIndex[10:0] ? 30'h3f5f5a5d : _GEN_1715; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1717 = 11'h2b4 == io_sinIndex[10:0] ? 30'h3f5f8b6f : _GEN_1716; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1718 = 11'h2b5 == io_sinIndex[10:0] ? 30'h3f5fbc5e : _GEN_1717; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1719 = 11'h2b6 == io_sinIndex[10:0] ? 30'h3f5fed2b : _GEN_1718; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1720 = 11'h2b7 == io_sinIndex[10:0] ? 30'h3f601dd6 : _GEN_1719; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1721 = 11'h2b8 == io_sinIndex[10:0] ? 30'h3f604e5e : _GEN_1720; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1722 = 11'h2b9 == io_sinIndex[10:0] ? 30'h3f607ec3 : _GEN_1721; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1723 = 11'h2ba == io_sinIndex[10:0] ? 30'h3f60af06 : _GEN_1722; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1724 = 11'h2bb == io_sinIndex[10:0] ? 30'h3f60df26 : _GEN_1723; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1725 = 11'h2bc == io_sinIndex[10:0] ? 30'h3f610f23 : _GEN_1724; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1726 = 11'h2bd == io_sinIndex[10:0] ? 30'h3f613efe : _GEN_1725; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1727 = 11'h2be == io_sinIndex[10:0] ? 30'h3f616eb5 : _GEN_1726; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1728 = 11'h2bf == io_sinIndex[10:0] ? 30'h3f619e4a : _GEN_1727; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1729 = 11'h2c0 == io_sinIndex[10:0] ? 30'h3f61cdbd : _GEN_1728; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1730 = 11'h2c1 == io_sinIndex[10:0] ? 30'h3f61fd0c : _GEN_1729; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1731 = 11'h2c2 == io_sinIndex[10:0] ? 30'h3f622c39 : _GEN_1730; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1732 = 11'h2c3 == io_sinIndex[10:0] ? 30'h3f625b42 : _GEN_1731; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1733 = 11'h2c4 == io_sinIndex[10:0] ? 30'h3f628a29 : _GEN_1732; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1734 = 11'h2c5 == io_sinIndex[10:0] ? 30'h3f62b8ed : _GEN_1733; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1735 = 11'h2c6 == io_sinIndex[10:0] ? 30'h3f62e78d : _GEN_1734; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1736 = 11'h2c7 == io_sinIndex[10:0] ? 30'h3f63160b : _GEN_1735; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1737 = 11'h2c8 == io_sinIndex[10:0] ? 30'h3f634466 : _GEN_1736; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1738 = 11'h2c9 == io_sinIndex[10:0] ? 30'h3f63729e : _GEN_1737; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1739 = 11'h2ca == io_sinIndex[10:0] ? 30'h3f63a0b2 : _GEN_1738; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1740 = 11'h2cb == io_sinIndex[10:0] ? 30'h3f63cea4 : _GEN_1739; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1741 = 11'h2cc == io_sinIndex[10:0] ? 30'h3f63fc72 : _GEN_1740; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1742 = 11'h2cd == io_sinIndex[10:0] ? 30'h3f642a1d : _GEN_1741; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1743 = 11'h2ce == io_sinIndex[10:0] ? 30'h3f6457a5 : _GEN_1742; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1744 = 11'h2cf == io_sinIndex[10:0] ? 30'h3f64850a : _GEN_1743; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1745 = 11'h2d0 == io_sinIndex[10:0] ? 30'h3f64b24b : _GEN_1744; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1746 = 11'h2d1 == io_sinIndex[10:0] ? 30'h3f64df69 : _GEN_1745; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1747 = 11'h2d2 == io_sinIndex[10:0] ? 30'h3f650c64 : _GEN_1746; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1748 = 11'h2d3 == io_sinIndex[10:0] ? 30'h3f65393b : _GEN_1747; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1749 = 11'h2d4 == io_sinIndex[10:0] ? 30'h3f6565f0 : _GEN_1748; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1750 = 11'h2d5 == io_sinIndex[10:0] ? 30'h3f659280 : _GEN_1749; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1751 = 11'h2d6 == io_sinIndex[10:0] ? 30'h3f65beee : _GEN_1750; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1752 = 11'h2d7 == io_sinIndex[10:0] ? 30'h3f65eb37 : _GEN_1751; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1753 = 11'h2d8 == io_sinIndex[10:0] ? 30'h3f66175e : _GEN_1752; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1754 = 11'h2d9 == io_sinIndex[10:0] ? 30'h3f664361 : _GEN_1753; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1755 = 11'h2da == io_sinIndex[10:0] ? 30'h3f666f40 : _GEN_1754; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1756 = 11'h2db == io_sinIndex[10:0] ? 30'h3f669afc : _GEN_1755; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1757 = 11'h2dc == io_sinIndex[10:0] ? 30'h3f66c694 : _GEN_1756; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1758 = 11'h2dd == io_sinIndex[10:0] ? 30'h3f66f209 : _GEN_1757; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1759 = 11'h2de == io_sinIndex[10:0] ? 30'h3f671d5a : _GEN_1758; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1760 = 11'h2df == io_sinIndex[10:0] ? 30'h3f674887 : _GEN_1759; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1761 = 11'h2e0 == io_sinIndex[10:0] ? 30'h3f677391 : _GEN_1760; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1762 = 11'h2e1 == io_sinIndex[10:0] ? 30'h3f679e77 : _GEN_1761; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1763 = 11'h2e2 == io_sinIndex[10:0] ? 30'h3f67c939 : _GEN_1762; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1764 = 11'h2e3 == io_sinIndex[10:0] ? 30'h3f67f3d7 : _GEN_1763; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1765 = 11'h2e4 == io_sinIndex[10:0] ? 30'h3f681e52 : _GEN_1764; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1766 = 11'h2e5 == io_sinIndex[10:0] ? 30'h3f6848a9 : _GEN_1765; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1767 = 11'h2e6 == io_sinIndex[10:0] ? 30'h3f6872dc : _GEN_1766; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1768 = 11'h2e7 == io_sinIndex[10:0] ? 30'h3f689ceb : _GEN_1767; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1769 = 11'h2e8 == io_sinIndex[10:0] ? 30'h3f68c6d6 : _GEN_1768; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1770 = 11'h2e9 == io_sinIndex[10:0] ? 30'h3f68f09e : _GEN_1769; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1771 = 11'h2ea == io_sinIndex[10:0] ? 30'h3f691a41 : _GEN_1770; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1772 = 11'h2eb == io_sinIndex[10:0] ? 30'h3f6943c0 : _GEN_1771; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1773 = 11'h2ec == io_sinIndex[10:0] ? 30'h3f696d1c : _GEN_1772; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1774 = 11'h2ed == io_sinIndex[10:0] ? 30'h3f699653 : _GEN_1773; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1775 = 11'h2ee == io_sinIndex[10:0] ? 30'h3f69bf67 : _GEN_1774; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1776 = 11'h2ef == io_sinIndex[10:0] ? 30'h3f69e856 : _GEN_1775; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1777 = 11'h2f0 == io_sinIndex[10:0] ? 30'h3f6a1121 : _GEN_1776; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1778 = 11'h2f1 == io_sinIndex[10:0] ? 30'h3f6a39c8 : _GEN_1777; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1779 = 11'h2f2 == io_sinIndex[10:0] ? 30'h3f6a624b : _GEN_1778; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1780 = 11'h2f3 == io_sinIndex[10:0] ? 30'h3f6a8aaa : _GEN_1779; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1781 = 11'h2f4 == io_sinIndex[10:0] ? 30'h3f6ab2e5 : _GEN_1780; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1782 = 11'h2f5 == io_sinIndex[10:0] ? 30'h3f6adafb : _GEN_1781; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1783 = 11'h2f6 == io_sinIndex[10:0] ? 30'h3f6b02ed : _GEN_1782; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1784 = 11'h2f7 == io_sinIndex[10:0] ? 30'h3f6b2abb : _GEN_1783; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1785 = 11'h2f8 == io_sinIndex[10:0] ? 30'h3f6b5265 : _GEN_1784; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1786 = 11'h2f9 == io_sinIndex[10:0] ? 30'h3f6b79ea : _GEN_1785; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1787 = 11'h2fa == io_sinIndex[10:0] ? 30'h3f6ba14b : _GEN_1786; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1788 = 11'h2fb == io_sinIndex[10:0] ? 30'h3f6bc888 : _GEN_1787; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1789 = 11'h2fc == io_sinIndex[10:0] ? 30'h3f6befa0 : _GEN_1788; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1790 = 11'h2fd == io_sinIndex[10:0] ? 30'h3f6c1694 : _GEN_1789; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1791 = 11'h2fe == io_sinIndex[10:0] ? 30'h3f6c3d63 : _GEN_1790; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1792 = 11'h2ff == io_sinIndex[10:0] ? 30'h3f6c640e : _GEN_1791; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1793 = 11'h300 == io_sinIndex[10:0] ? 30'h3f6c8a95 : _GEN_1792; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1794 = 11'h301 == io_sinIndex[10:0] ? 30'h3f6cb0f7 : _GEN_1793; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1795 = 11'h302 == io_sinIndex[10:0] ? 30'h3f6cd734 : _GEN_1794; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1796 = 11'h303 == io_sinIndex[10:0] ? 30'h3f6cfd4d : _GEN_1795; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1797 = 11'h304 == io_sinIndex[10:0] ? 30'h3f6d2342 : _GEN_1796; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1798 = 11'h305 == io_sinIndex[10:0] ? 30'h3f6d4912 : _GEN_1797; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1799 = 11'h306 == io_sinIndex[10:0] ? 30'h3f6d6ebd : _GEN_1798; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1800 = 11'h307 == io_sinIndex[10:0] ? 30'h3f6d9443 : _GEN_1799; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1801 = 11'h308 == io_sinIndex[10:0] ? 30'h3f6db9a5 : _GEN_1800; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1802 = 11'h309 == io_sinIndex[10:0] ? 30'h3f6ddee3 : _GEN_1801; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1803 = 11'h30a == io_sinIndex[10:0] ? 30'h3f6e03fb : _GEN_1802; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1804 = 11'h30b == io_sinIndex[10:0] ? 30'h3f6e28ef : _GEN_1803; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1805 = 11'h30c == io_sinIndex[10:0] ? 30'h3f6e4dbe : _GEN_1804; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1806 = 11'h30d == io_sinIndex[10:0] ? 30'h3f6e7268 : _GEN_1805; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1807 = 11'h30e == io_sinIndex[10:0] ? 30'h3f6e96ee : _GEN_1806; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1808 = 11'h30f == io_sinIndex[10:0] ? 30'h3f6ebb4e : _GEN_1807; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1809 = 11'h310 == io_sinIndex[10:0] ? 30'h3f6edf8a : _GEN_1808; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1810 = 11'h311 == io_sinIndex[10:0] ? 30'h3f6f03a1 : _GEN_1809; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1811 = 11'h312 == io_sinIndex[10:0] ? 30'h3f6f2793 : _GEN_1810; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1812 = 11'h313 == io_sinIndex[10:0] ? 30'h3f6f4b61 : _GEN_1811; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1813 = 11'h314 == io_sinIndex[10:0] ? 30'h3f6f6f09 : _GEN_1812; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1814 = 11'h315 == io_sinIndex[10:0] ? 30'h3f6f928c : _GEN_1813; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1815 = 11'h316 == io_sinIndex[10:0] ? 30'h3f6fb5eb : _GEN_1814; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1816 = 11'h317 == io_sinIndex[10:0] ? 30'h3f6fd924 : _GEN_1815; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1817 = 11'h318 == io_sinIndex[10:0] ? 30'h3f6ffc39 : _GEN_1816; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1818 = 11'h319 == io_sinIndex[10:0] ? 30'h3f701f28 : _GEN_1817; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1819 = 11'h31a == io_sinIndex[10:0] ? 30'h3f7041f2 : _GEN_1818; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1820 = 11'h31b == io_sinIndex[10:0] ? 30'h3f706498 : _GEN_1819; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1821 = 11'h31c == io_sinIndex[10:0] ? 30'h3f708718 : _GEN_1820; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1822 = 11'h31d == io_sinIndex[10:0] ? 30'h3f70a973 : _GEN_1821; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1823 = 11'h31e == io_sinIndex[10:0] ? 30'h3f70cba9 : _GEN_1822; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1824 = 11'h31f == io_sinIndex[10:0] ? 30'h3f70edba : _GEN_1823; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1825 = 11'h320 == io_sinIndex[10:0] ? 30'h3f710fa5 : _GEN_1824; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1826 = 11'h321 == io_sinIndex[10:0] ? 30'h3f71316c : _GEN_1825; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1827 = 11'h322 == io_sinIndex[10:0] ? 30'h3f71530d : _GEN_1826; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1828 = 11'h323 == io_sinIndex[10:0] ? 30'h3f717489 : _GEN_1827; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1829 = 11'h324 == io_sinIndex[10:0] ? 30'h3f7195e0 : _GEN_1828; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1830 = 11'h325 == io_sinIndex[10:0] ? 30'h3f71b711 : _GEN_1829; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1831 = 11'h326 == io_sinIndex[10:0] ? 30'h3f71d81d : _GEN_1830; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1832 = 11'h327 == io_sinIndex[10:0] ? 30'h3f71f904 : _GEN_1831; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1833 = 11'h328 == io_sinIndex[10:0] ? 30'h3f7219c6 : _GEN_1832; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1834 = 11'h329 == io_sinIndex[10:0] ? 30'h3f723a62 : _GEN_1833; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1835 = 11'h32a == io_sinIndex[10:0] ? 30'h3f725ad9 : _GEN_1834; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1836 = 11'h32b == io_sinIndex[10:0] ? 30'h3f727b2a : _GEN_1835; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1837 = 11'h32c == io_sinIndex[10:0] ? 30'h3f729b56 : _GEN_1836; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1838 = 11'h32d == io_sinIndex[10:0] ? 30'h3f72bb5c : _GEN_1837; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1839 = 11'h32e == io_sinIndex[10:0] ? 30'h3f72db3e : _GEN_1838; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1840 = 11'h32f == io_sinIndex[10:0] ? 30'h3f72faf9 : _GEN_1839; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1841 = 11'h330 == io_sinIndex[10:0] ? 30'h3f731a8f : _GEN_1840; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1842 = 11'h331 == io_sinIndex[10:0] ? 30'h3f733a00 : _GEN_1841; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1843 = 11'h332 == io_sinIndex[10:0] ? 30'h3f73594b : _GEN_1842; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1844 = 11'h333 == io_sinIndex[10:0] ? 30'h3f737871 : _GEN_1843; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1845 = 11'h334 == io_sinIndex[10:0] ? 30'h3f739771 : _GEN_1844; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1846 = 11'h335 == io_sinIndex[10:0] ? 30'h3f73b64b : _GEN_1845; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1847 = 11'h336 == io_sinIndex[10:0] ? 30'h3f73d500 : _GEN_1846; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1848 = 11'h337 == io_sinIndex[10:0] ? 30'h3f73f38f : _GEN_1847; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1849 = 11'h338 == io_sinIndex[10:0] ? 30'h3f7411f9 : _GEN_1848; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1850 = 11'h339 == io_sinIndex[10:0] ? 30'h3f74303c : _GEN_1849; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1851 = 11'h33a == io_sinIndex[10:0] ? 30'h3f744e5b : _GEN_1850; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1852 = 11'h33b == io_sinIndex[10:0] ? 30'h3f746c53 : _GEN_1851; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1853 = 11'h33c == io_sinIndex[10:0] ? 30'h3f748a26 : _GEN_1852; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1854 = 11'h33d == io_sinIndex[10:0] ? 30'h3f74a7d3 : _GEN_1853; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1855 = 11'h33e == io_sinIndex[10:0] ? 30'h3f74c55a : _GEN_1854; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1856 = 11'h33f == io_sinIndex[10:0] ? 30'h3f74e2bc : _GEN_1855; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1857 = 11'h340 == io_sinIndex[10:0] ? 30'h3f74fff8 : _GEN_1856; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1858 = 11'h341 == io_sinIndex[10:0] ? 30'h3f751d0e : _GEN_1857; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1859 = 11'h342 == io_sinIndex[10:0] ? 30'h3f7539fe : _GEN_1858; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1860 = 11'h343 == io_sinIndex[10:0] ? 30'h3f7556c8 : _GEN_1859; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1861 = 11'h344 == io_sinIndex[10:0] ? 30'h3f75736d : _GEN_1860; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1862 = 11'h345 == io_sinIndex[10:0] ? 30'h3f758feb : _GEN_1861; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1863 = 11'h346 == io_sinIndex[10:0] ? 30'h3f75ac44 : _GEN_1862; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1864 = 11'h347 == io_sinIndex[10:0] ? 30'h3f75c877 : _GEN_1863; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1865 = 11'h348 == io_sinIndex[10:0] ? 30'h3f75e484 : _GEN_1864; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1866 = 11'h349 == io_sinIndex[10:0] ? 30'h3f76006b : _GEN_1865; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1867 = 11'h34a == io_sinIndex[10:0] ? 30'h3f761c2c : _GEN_1866; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1868 = 11'h34b == io_sinIndex[10:0] ? 30'h3f7637c7 : _GEN_1867; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1869 = 11'h34c == io_sinIndex[10:0] ? 30'h3f76533c : _GEN_1868; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1870 = 11'h34d == io_sinIndex[10:0] ? 30'h3f766e8b : _GEN_1869; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1871 = 11'h34e == io_sinIndex[10:0] ? 30'h3f7689b4 : _GEN_1870; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1872 = 11'h34f == io_sinIndex[10:0] ? 30'h3f76a4b7 : _GEN_1871; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1873 = 11'h350 == io_sinIndex[10:0] ? 30'h3f76bf94 : _GEN_1872; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1874 = 11'h351 == io_sinIndex[10:0] ? 30'h3f76da4b : _GEN_1873; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1875 = 11'h352 == io_sinIndex[10:0] ? 30'h3f76f4db : _GEN_1874; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1876 = 11'h353 == io_sinIndex[10:0] ? 30'h3f770f46 : _GEN_1875; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1877 = 11'h354 == io_sinIndex[10:0] ? 30'h3f77298b : _GEN_1876; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1878 = 11'h355 == io_sinIndex[10:0] ? 30'h3f7743a9 : _GEN_1877; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1879 = 11'h356 == io_sinIndex[10:0] ? 30'h3f775da1 : _GEN_1878; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1880 = 11'h357 == io_sinIndex[10:0] ? 30'h3f777773 : _GEN_1879; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1881 = 11'h358 == io_sinIndex[10:0] ? 30'h3f77911f : _GEN_1880; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1882 = 11'h359 == io_sinIndex[10:0] ? 30'h3f77aaa5 : _GEN_1881; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1883 = 11'h35a == io_sinIndex[10:0] ? 30'h3f77c405 : _GEN_1882; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1884 = 11'h35b == io_sinIndex[10:0] ? 30'h3f77dd3e : _GEN_1883; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1885 = 11'h35c == io_sinIndex[10:0] ? 30'h3f77f651 : _GEN_1884; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1886 = 11'h35d == io_sinIndex[10:0] ? 30'h3f780f3e : _GEN_1885; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1887 = 11'h35e == io_sinIndex[10:0] ? 30'h3f782804 : _GEN_1886; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1888 = 11'h35f == io_sinIndex[10:0] ? 30'h3f7840a4 : _GEN_1887; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1889 = 11'h360 == io_sinIndex[10:0] ? 30'h3f78591e : _GEN_1888; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1890 = 11'h361 == io_sinIndex[10:0] ? 30'h3f787172 : _GEN_1889; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1891 = 11'h362 == io_sinIndex[10:0] ? 30'h3f78899f : _GEN_1890; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1892 = 11'h363 == io_sinIndex[10:0] ? 30'h3f78a1a6 : _GEN_1891; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1893 = 11'h364 == io_sinIndex[10:0] ? 30'h3f78b987 : _GEN_1892; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1894 = 11'h365 == io_sinIndex[10:0] ? 30'h3f78d141 : _GEN_1893; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1895 = 11'h366 == io_sinIndex[10:0] ? 30'h3f78e8d5 : _GEN_1894; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1896 = 11'h367 == io_sinIndex[10:0] ? 30'h3f790042 : _GEN_1895; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1897 = 11'h368 == io_sinIndex[10:0] ? 30'h3f791789 : _GEN_1896; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1898 = 11'h369 == io_sinIndex[10:0] ? 30'h3f792eaa : _GEN_1897; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1899 = 11'h36a == io_sinIndex[10:0] ? 30'h3f7945a4 : _GEN_1898; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1900 = 11'h36b == io_sinIndex[10:0] ? 30'h3f795c77 : _GEN_1899; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1901 = 11'h36c == io_sinIndex[10:0] ? 30'h3f797325 : _GEN_1900; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1902 = 11'h36d == io_sinIndex[10:0] ? 30'h3f7989ab : _GEN_1901; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1903 = 11'h36e == io_sinIndex[10:0] ? 30'h3f79a00b : _GEN_1902; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1904 = 11'h36f == io_sinIndex[10:0] ? 30'h3f79b645 : _GEN_1903; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1905 = 11'h370 == io_sinIndex[10:0] ? 30'h3f79cc58 : _GEN_1904; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1906 = 11'h371 == io_sinIndex[10:0] ? 30'h3f79e245 : _GEN_1905; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1907 = 11'h372 == io_sinIndex[10:0] ? 30'h3f79f80b : _GEN_1906; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1908 = 11'h373 == io_sinIndex[10:0] ? 30'h3f7a0daa : _GEN_1907; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1909 = 11'h374 == io_sinIndex[10:0] ? 30'h3f7a2323 : _GEN_1908; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1910 = 11'h375 == io_sinIndex[10:0] ? 30'h3f7a3876 : _GEN_1909; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1911 = 11'h376 == io_sinIndex[10:0] ? 30'h3f7a4da1 : _GEN_1910; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1912 = 11'h377 == io_sinIndex[10:0] ? 30'h3f7a62a6 : _GEN_1911; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1913 = 11'h378 == io_sinIndex[10:0] ? 30'h3f7a7785 : _GEN_1912; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1914 = 11'h379 == io_sinIndex[10:0] ? 30'h3f7a8c3d : _GEN_1913; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1915 = 11'h37a == io_sinIndex[10:0] ? 30'h3f7aa0ce : _GEN_1914; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1916 = 11'h37b == io_sinIndex[10:0] ? 30'h3f7ab538 : _GEN_1915; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1917 = 11'h37c == io_sinIndex[10:0] ? 30'h3f7ac97c : _GEN_1916; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1918 = 11'h37d == io_sinIndex[10:0] ? 30'h3f7add99 : _GEN_1917; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1919 = 11'h37e == io_sinIndex[10:0] ? 30'h3f7af190 : _GEN_1918; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1920 = 11'h37f == io_sinIndex[10:0] ? 30'h3f7b055f : _GEN_1919; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1921 = 11'h380 == io_sinIndex[10:0] ? 30'h3f7b1908 : _GEN_1920; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1922 = 11'h381 == io_sinIndex[10:0] ? 30'h3f7b2c8a : _GEN_1921; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1923 = 11'h382 == io_sinIndex[10:0] ? 30'h3f7b3fe6 : _GEN_1922; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1924 = 11'h383 == io_sinIndex[10:0] ? 30'h3f7b531b : _GEN_1923; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1925 = 11'h384 == io_sinIndex[10:0] ? 30'h3f7b6628 : _GEN_1924; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1926 = 11'h385 == io_sinIndex[10:0] ? 30'h3f7b7910 : _GEN_1925; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1927 = 11'h386 == io_sinIndex[10:0] ? 30'h3f7b8bd0 : _GEN_1926; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1928 = 11'h387 == io_sinIndex[10:0] ? 30'h3f7b9e69 : _GEN_1927; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1929 = 11'h388 == io_sinIndex[10:0] ? 30'h3f7bb0dc : _GEN_1928; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1930 = 11'h389 == io_sinIndex[10:0] ? 30'h3f7bc328 : _GEN_1929; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1931 = 11'h38a == io_sinIndex[10:0] ? 30'h3f7bd54d : _GEN_1930; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1932 = 11'h38b == io_sinIndex[10:0] ? 30'h3f7be74b : _GEN_1931; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1933 = 11'h38c == io_sinIndex[10:0] ? 30'h3f7bf922 : _GEN_1932; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1934 = 11'h38d == io_sinIndex[10:0] ? 30'h3f7c0ad3 : _GEN_1933; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1935 = 11'h38e == io_sinIndex[10:0] ? 30'h3f7c1c5c : _GEN_1934; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1936 = 11'h38f == io_sinIndex[10:0] ? 30'h3f7c2dbf : _GEN_1935; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1937 = 11'h390 == io_sinIndex[10:0] ? 30'h3f7c3efb : _GEN_1936; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1938 = 11'h391 == io_sinIndex[10:0] ? 30'h3f7c5010 : _GEN_1937; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1939 = 11'h392 == io_sinIndex[10:0] ? 30'h3f7c60fd : _GEN_1938; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1940 = 11'h393 == io_sinIndex[10:0] ? 30'h3f7c71c4 : _GEN_1939; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1941 = 11'h394 == io_sinIndex[10:0] ? 30'h3f7c8264 : _GEN_1940; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1942 = 11'h395 == io_sinIndex[10:0] ? 30'h3f7c92dd : _GEN_1941; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1943 = 11'h396 == io_sinIndex[10:0] ? 30'h3f7ca32f : _GEN_1942; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1944 = 11'h397 == io_sinIndex[10:0] ? 30'h3f7cb35b : _GEN_1943; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1945 = 11'h398 == io_sinIndex[10:0] ? 30'h3f7cc35f : _GEN_1944; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1946 = 11'h399 == io_sinIndex[10:0] ? 30'h3f7cd33c : _GEN_1945; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1947 = 11'h39a == io_sinIndex[10:0] ? 30'h3f7ce2f2 : _GEN_1946; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1948 = 11'h39b == io_sinIndex[10:0] ? 30'h3f7cf281 : _GEN_1947; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1949 = 11'h39c == io_sinIndex[10:0] ? 30'h3f7d01e9 : _GEN_1948; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1950 = 11'h39d == io_sinIndex[10:0] ? 30'h3f7d112a : _GEN_1949; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1951 = 11'h39e == io_sinIndex[10:0] ? 30'h3f7d2044 : _GEN_1950; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1952 = 11'h39f == io_sinIndex[10:0] ? 30'h3f7d2f37 : _GEN_1951; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1953 = 11'h3a0 == io_sinIndex[10:0] ? 30'h3f7d3e03 : _GEN_1952; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1954 = 11'h3a1 == io_sinIndex[10:0] ? 30'h3f7d4ca8 : _GEN_1953; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1955 = 11'h3a2 == io_sinIndex[10:0] ? 30'h3f7d5b25 : _GEN_1954; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1956 = 11'h3a3 == io_sinIndex[10:0] ? 30'h3f7d697c : _GEN_1955; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1957 = 11'h3a4 == io_sinIndex[10:0] ? 30'h3f7d77ab : _GEN_1956; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1958 = 11'h3a5 == io_sinIndex[10:0] ? 30'h3f7d85b4 : _GEN_1957; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1959 = 11'h3a6 == io_sinIndex[10:0] ? 30'h3f7d9395 : _GEN_1958; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1960 = 11'h3a7 == io_sinIndex[10:0] ? 30'h3f7da14f : _GEN_1959; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1961 = 11'h3a8 == io_sinIndex[10:0] ? 30'h3f7daee2 : _GEN_1960; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1962 = 11'h3a9 == io_sinIndex[10:0] ? 30'h3f7dbc4e : _GEN_1961; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1963 = 11'h3aa == io_sinIndex[10:0] ? 30'h3f7dc993 : _GEN_1962; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1964 = 11'h3ab == io_sinIndex[10:0] ? 30'h3f7dd6b0 : _GEN_1963; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1965 = 11'h3ac == io_sinIndex[10:0] ? 30'h3f7de3a7 : _GEN_1964; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1966 = 11'h3ad == io_sinIndex[10:0] ? 30'h3f7df076 : _GEN_1965; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1967 = 11'h3ae == io_sinIndex[10:0] ? 30'h3f7dfd1e : _GEN_1966; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1968 = 11'h3af == io_sinIndex[10:0] ? 30'h3f7e099f : _GEN_1967; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1969 = 11'h3b0 == io_sinIndex[10:0] ? 30'h3f7e15f9 : _GEN_1968; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1970 = 11'h3b1 == io_sinIndex[10:0] ? 30'h3f7e222b : _GEN_1969; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1971 = 11'h3b2 == io_sinIndex[10:0] ? 30'h3f7e2e36 : _GEN_1970; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1972 = 11'h3b3 == io_sinIndex[10:0] ? 30'h3f7e3a1b : _GEN_1971; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1973 = 11'h3b4 == io_sinIndex[10:0] ? 30'h3f7e45d7 : _GEN_1972; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1974 = 11'h3b5 == io_sinIndex[10:0] ? 30'h3f7e516d : _GEN_1973; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1975 = 11'h3b6 == io_sinIndex[10:0] ? 30'h3f7e5cdb : _GEN_1974; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1976 = 11'h3b7 == io_sinIndex[10:0] ? 30'h3f7e6822 : _GEN_1975; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1977 = 11'h3b8 == io_sinIndex[10:0] ? 30'h3f7e7342 : _GEN_1976; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1978 = 11'h3b9 == io_sinIndex[10:0] ? 30'h3f7e7e3b : _GEN_1977; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1979 = 11'h3ba == io_sinIndex[10:0] ? 30'h3f7e890c : _GEN_1978; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1980 = 11'h3bb == io_sinIndex[10:0] ? 30'h3f7e93b6 : _GEN_1979; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1981 = 11'h3bc == io_sinIndex[10:0] ? 30'h3f7e9e39 : _GEN_1980; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1982 = 11'h3bd == io_sinIndex[10:0] ? 30'h3f7ea895 : _GEN_1981; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1983 = 11'h3be == io_sinIndex[10:0] ? 30'h3f7eb2c9 : _GEN_1982; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1984 = 11'h3bf == io_sinIndex[10:0] ? 30'h3f7ebcd6 : _GEN_1983; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1985 = 11'h3c0 == io_sinIndex[10:0] ? 30'h3f7ec6bb : _GEN_1984; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1986 = 11'h3c1 == io_sinIndex[10:0] ? 30'h3f7ed07a : _GEN_1985; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1987 = 11'h3c2 == io_sinIndex[10:0] ? 30'h3f7eda11 : _GEN_1986; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1988 = 11'h3c3 == io_sinIndex[10:0] ? 30'h3f7ee380 : _GEN_1987; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1989 = 11'h3c4 == io_sinIndex[10:0] ? 30'h3f7eecc9 : _GEN_1988; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1990 = 11'h3c5 == io_sinIndex[10:0] ? 30'h3f7ef5ea : _GEN_1989; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1991 = 11'h3c6 == io_sinIndex[10:0] ? 30'h3f7efee3 : _GEN_1990; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1992 = 11'h3c7 == io_sinIndex[10:0] ? 30'h3f7f07b6 : _GEN_1991; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1993 = 11'h3c8 == io_sinIndex[10:0] ? 30'h3f7f1061 : _GEN_1992; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1994 = 11'h3c9 == io_sinIndex[10:0] ? 30'h3f7f18e4 : _GEN_1993; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1995 = 11'h3ca == io_sinIndex[10:0] ? 30'h3f7f2141 : _GEN_1994; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1996 = 11'h3cb == io_sinIndex[10:0] ? 30'h3f7f2976 : _GEN_1995; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1997 = 11'h3cc == io_sinIndex[10:0] ? 30'h3f7f3183 : _GEN_1996; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1998 = 11'h3cd == io_sinIndex[10:0] ? 30'h3f7f3969 : _GEN_1997; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_1999 = 11'h3ce == io_sinIndex[10:0] ? 30'h3f7f4128 : _GEN_1998; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2000 = 11'h3cf == io_sinIndex[10:0] ? 30'h3f7f48c0 : _GEN_1999; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2001 = 11'h3d0 == io_sinIndex[10:0] ? 30'h3f7f5030 : _GEN_2000; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2002 = 11'h3d1 == io_sinIndex[10:0] ? 30'h3f7f5778 : _GEN_2001; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2003 = 11'h3d2 == io_sinIndex[10:0] ? 30'h3f7f5e99 : _GEN_2002; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2004 = 11'h3d3 == io_sinIndex[10:0] ? 30'h3f7f6593 : _GEN_2003; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2005 = 11'h3d4 == io_sinIndex[10:0] ? 30'h3f7f6c66 : _GEN_2004; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2006 = 11'h3d5 == io_sinIndex[10:0] ? 30'h3f7f7311 : _GEN_2005; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2007 = 11'h3d6 == io_sinIndex[10:0] ? 30'h3f7f7994 : _GEN_2006; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2008 = 11'h3d7 == io_sinIndex[10:0] ? 30'h3f7f7ff0 : _GEN_2007; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2009 = 11'h3d8 == io_sinIndex[10:0] ? 30'h3f7f8625 : _GEN_2008; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2010 = 11'h3d9 == io_sinIndex[10:0] ? 30'h3f7f8c33 : _GEN_2009; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2011 = 11'h3da == io_sinIndex[10:0] ? 30'h3f7f9219 : _GEN_2010; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2012 = 11'h3db == io_sinIndex[10:0] ? 30'h3f7f97d7 : _GEN_2011; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2013 = 11'h3dc == io_sinIndex[10:0] ? 30'h3f7f9d6e : _GEN_2012; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2014 = 11'h3dd == io_sinIndex[10:0] ? 30'h3f7fa2de : _GEN_2013; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2015 = 11'h3de == io_sinIndex[10:0] ? 30'h3f7fa826 : _GEN_2014; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2016 = 11'h3df == io_sinIndex[10:0] ? 30'h3f7fad47 : _GEN_2015; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2017 = 11'h3e0 == io_sinIndex[10:0] ? 30'h3f7fb240 : _GEN_2016; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2018 = 11'h3e1 == io_sinIndex[10:0] ? 30'h3f7fb712 : _GEN_2017; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2019 = 11'h3e2 == io_sinIndex[10:0] ? 30'h3f7fbbbc : _GEN_2018; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2020 = 11'h3e3 == io_sinIndex[10:0] ? 30'h3f7fc03f : _GEN_2019; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2021 = 11'h3e4 == io_sinIndex[10:0] ? 30'h3f7fc49a : _GEN_2020; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2022 = 11'h3e5 == io_sinIndex[10:0] ? 30'h3f7fc8ce : _GEN_2021; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2023 = 11'h3e6 == io_sinIndex[10:0] ? 30'h3f7fccdb : _GEN_2022; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2024 = 11'h3e7 == io_sinIndex[10:0] ? 30'h3f7fd0c0 : _GEN_2023; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2025 = 11'h3e8 == io_sinIndex[10:0] ? 30'h3f7fd47e : _GEN_2024; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2026 = 11'h3e9 == io_sinIndex[10:0] ? 30'h3f7fd814 : _GEN_2025; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2027 = 11'h3ea == io_sinIndex[10:0] ? 30'h3f7fdb82 : _GEN_2026; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2028 = 11'h3eb == io_sinIndex[10:0] ? 30'h3f7fdeca : _GEN_2027; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2029 = 11'h3ec == io_sinIndex[10:0] ? 30'h3f7fe1e9 : _GEN_2028; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2030 = 11'h3ed == io_sinIndex[10:0] ? 30'h3f7fe4e2 : _GEN_2029; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2031 = 11'h3ee == io_sinIndex[10:0] ? 30'h3f7fe7b2 : _GEN_2030; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2032 = 11'h3ef == io_sinIndex[10:0] ? 30'h3f7fea5c : _GEN_2031; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2033 = 11'h3f0 == io_sinIndex[10:0] ? 30'h3f7fecdd : _GEN_2032; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2034 = 11'h3f1 == io_sinIndex[10:0] ? 30'h3f7fef38 : _GEN_2033; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2035 = 11'h3f2 == io_sinIndex[10:0] ? 30'h3f7ff16a : _GEN_2034; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2036 = 11'h3f3 == io_sinIndex[10:0] ? 30'h3f7ff376 : _GEN_2035; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2037 = 11'h3f4 == io_sinIndex[10:0] ? 30'h3f7ff559 : _GEN_2036; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2038 = 11'h3f5 == io_sinIndex[10:0] ? 30'h3f7ff716 : _GEN_2037; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2039 = 11'h3f6 == io_sinIndex[10:0] ? 30'h3f7ff8ab : _GEN_2038; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2040 = 11'h3f7 == io_sinIndex[10:0] ? 30'h3f7ffa18 : _GEN_2039; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2041 = 11'h3f8 == io_sinIndex[10:0] ? 30'h3f7ffb5e : _GEN_2040; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2042 = 11'h3f9 == io_sinIndex[10:0] ? 30'h3f7ffc7c : _GEN_2041; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2043 = 11'h3fa == io_sinIndex[10:0] ? 30'h3f7ffd73 : _GEN_2042; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2044 = 11'h3fb == io_sinIndex[10:0] ? 30'h3f7ffe42 : _GEN_2043; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2045 = 11'h3fc == io_sinIndex[10:0] ? 30'h3f7ffeea : _GEN_2044; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2046 = 11'h3fd == io_sinIndex[10:0] ? 30'h3f7fff6b : _GEN_2045; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2047 = 11'h3fe == io_sinIndex[10:0] ? 30'h3f7fffc4 : _GEN_2046; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2048 = 11'h3ff == io_sinIndex[10:0] ? 30'h3f7ffff5 : _GEN_2047; // @[LUTbank.scala 294:{21,21}]
  wire [29:0] _GEN_2049 = 11'h400 == io_sinIndex[10:0] ? 30'h3f800000 : _GEN_2048; // @[LUTbank.scala 294:{21,21}]
  assign io_sinOut = io_EN ? {{2'd0}, _GEN_2049} : 32'h0; // @[LUTbank.scala 294:21]
  assign io_cosOut = io_EN ? {{2'd0}, _GEN_1024} : 32'h0; // @[LUTbank.scala 293:21]
  assign io_ENout = io_EN; // @[LUTbank.scala 295:21]
endmodule
module SinCosLUT(
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_angle,
  output [31:0] io_sinOut,
  output [31:0] io_cosOut,
  output        io_ENout,
  output [31:0] io_xFWD_0,
  output [31:0] io_xFWD_1
);
  wire  indexCalculator_io_EN; // @[sincosLUT.scala 92:31]
  wire [31:0] indexCalculator_io_angle; // @[sincosLUT.scala 92:31]
  wire [31:0] indexCalculator_io_cosIndex; // @[sincosLUT.scala 92:31]
  wire [31:0] indexCalculator_io_sinIndex; // @[sincosLUT.scala 92:31]
  wire  indexCalculator_io_cosSign; // @[sincosLUT.scala 92:31]
  wire  indexCalculator_io_sinSign; // @[sincosLUT.scala 92:31]
  wire  indexCalculator_io_ENout; // @[sincosLUT.scala 92:31]
  wire  lutModule_io_EN; // @[sincosLUT.scala 93:25]
  wire [31:0] lutModule_io_cosIndex; // @[sincosLUT.scala 93:25]
  wire [31:0] lutModule_io_sinIndex; // @[sincosLUT.scala 93:25]
  wire [31:0] lutModule_io_sinOut; // @[sincosLUT.scala 93:25]
  wire [31:0] lutModule_io_cosOut; // @[sincosLUT.scala 93:25]
  wire  lutModule_io_ENout; // @[sincosLUT.scala 93:25]
  wire [31:0] _io_cosOut_T_1 = {indexCalculator_io_cosSign,lutModule_io_cosOut[30:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_sinOut_T_1 = {indexCalculator_io_sinSign,lutModule_io_sinOut[30:0]}; // @[Cat.scala 33:92]
  IndexCalculator indexCalculator ( // @[sincosLUT.scala 92:31]
    .io_EN(indexCalculator_io_EN),
    .io_angle(indexCalculator_io_angle),
    .io_cosIndex(indexCalculator_io_cosIndex),
    .io_sinIndex(indexCalculator_io_sinIndex),
    .io_cosSign(indexCalculator_io_cosSign),
    .io_sinSign(indexCalculator_io_sinSign),
    .io_ENout(indexCalculator_io_ENout)
  );
  CosLUT lutModule ( // @[sincosLUT.scala 93:25]
    .io_EN(lutModule_io_EN),
    .io_cosIndex(lutModule_io_cosIndex),
    .io_sinIndex(lutModule_io_sinIndex),
    .io_sinOut(lutModule_io_sinOut),
    .io_cosOut(lutModule_io_cosOut),
    .io_ENout(lutModule_io_ENout)
  );
  assign io_sinOut = lutModule_io_ENout ? _io_sinOut_T_1 : 32'h0; // @[sincosLUT.scala 106:19]
  assign io_cosOut = lutModule_io_ENout ? _io_cosOut_T_1 : 32'h0; // @[sincosLUT.scala 105:19]
  assign io_ENout = lutModule_io_ENout; // @[sincosLUT.scala 107:19]
  assign io_xFWD_0 = lutModule_io_ENout ? io_x_0 : 32'h0; // @[sincosLUT.scala 102:20]
  assign io_xFWD_1 = lutModule_io_ENout ? io_x_1 : 32'h0; // @[sincosLUT.scala 103:20]
  assign indexCalculator_io_EN = io_EN; // @[sincosLUT.scala 95:25]
  assign indexCalculator_io_angle = io_angle; // @[sincosLUT.scala 96:28]
  assign lutModule_io_EN = indexCalculator_io_ENout; // @[sincosLUT.scala 100:19]
  assign lutModule_io_cosIndex = indexCalculator_io_cosIndex; // @[sincosLUT.scala 98:25]
  assign lutModule_io_sinIndex = indexCalculator_io_sinIndex; // @[sincosLUT.scala 99:25]
endmodule
module FP32Adder(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire  adder_io_subOp; // @[FPU.scala 17:23]
  wire [32:0] adder_io_a; // @[FPU.scala 17:23]
  wire [32:0] adder_io_b; // @[FPU.scala 17:23]
  wire [32:0] adder_io_out; // @[FPU.scala 17:23]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = adder_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = adder_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,adder_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  AddRecFN adder ( // @[FPU.scala 17:23]
    .io_subOp(adder_io_subOp),
    .io_a(adder_io_a),
    .io_b(adder_io_b),
    .io_out(adder_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign adder_io_subOp = 1'h0; // @[FPU.scala 24:20]
  assign adder_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign adder_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module FP32RoPEcore(
  input         clock,
  input         reset,
  input         io_EN,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input  [31:0] io_sin,
  input  [31:0] io_cos,
  output [31:0] io_xhat_0,
  output [31:0] io_xhat_1,
  output        io_ENout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] FP32Mult0_io_a; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult0_io_b; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult0_io_result; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult1_io_a; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult1_io_b; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult1_io_result; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult2_io_a; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult2_io_b; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult2_io_result; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult3_io_a; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Mult3_io_b; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Mult3_io_result; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Sub_io_a; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32Sub_io_b; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32Sub_io_result; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32add_io_a; // @[RoPEModuleFP32.scala 135:25]
  wire [31:0] FP32add_io_b; // @[RoPEModuleFP32.scala 135:25]
  wire [31:0] FP32add_io_result; // @[RoPEModuleFP32.scala 135:25]
  reg [31:0] stage1Reg_0; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_1; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_2; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_3; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage2Reg_0; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_1; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_2; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_3; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage3Reg_0; // @[RoPEModuleFP32.scala 97:28]
  reg [31:0] stage3Reg_1; // @[RoPEModuleFP32.scala 97:28]
  reg  enReg_0; // @[RoPEModuleFP32.scala 98:24]
  reg  enReg_1; // @[RoPEModuleFP32.scala 98:24]
  reg  enReg_2; // @[RoPEModuleFP32.scala 98:24]
  wire [31:0] _WIRE_1_0 = FP32Sub_io_result; // @[RoPEModuleFP32.scala 139:{25,25}]
  wire [31:0] _WIRE_1_1 = FP32add_io_result; // @[RoPEModuleFP32.scala 139:{25,25}]
  FP32Multiplier FP32Mult0 ( // @[RoPEModuleFP32.scala 106:27]
    .io_a(FP32Mult0_io_a),
    .io_b(FP32Mult0_io_b),
    .io_result(FP32Mult0_io_result)
  );
  FP32Multiplier FP32Mult1 ( // @[RoPEModuleFP32.scala 110:27]
    .io_a(FP32Mult1_io_a),
    .io_b(FP32Mult1_io_b),
    .io_result(FP32Mult1_io_result)
  );
  FP32Multiplier FP32Mult2 ( // @[RoPEModuleFP32.scala 114:27]
    .io_a(FP32Mult2_io_a),
    .io_b(FP32Mult2_io_b),
    .io_result(FP32Mult2_io_result)
  );
  FP32Multiplier FP32Mult3 ( // @[RoPEModuleFP32.scala 118:27]
    .io_a(FP32Mult3_io_a),
    .io_b(FP32Mult3_io_b),
    .io_result(FP32Mult3_io_result)
  );
  FP32Sub FP32Sub ( // @[RoPEModuleFP32.scala 131:25]
    .io_a(FP32Sub_io_a),
    .io_b(FP32Sub_io_b),
    .io_result(FP32Sub_io_result)
  );
  FP32Adder FP32add ( // @[RoPEModuleFP32.scala 135:25]
    .io_a(FP32add_io_a),
    .io_b(FP32add_io_b),
    .io_result(FP32add_io_result)
  );
  assign io_xhat_0 = enReg_2 ? stage3Reg_0 : 32'h0; // @[RoPEModuleFP32.scala 142:22]
  assign io_xhat_1 = enReg_2 ? stage3Reg_1 : 32'h0; // @[RoPEModuleFP32.scala 143:22]
  assign io_ENout = enReg_2; // @[RoPEModuleFP32.scala 144:14]
  assign FP32Mult0_io_a = stage1Reg_0; // @[RoPEModuleFP32.scala 107:20]
  assign FP32Mult0_io_b = stage1Reg_2; // @[RoPEModuleFP32.scala 108:20]
  assign FP32Mult1_io_a = stage1Reg_1; // @[RoPEModuleFP32.scala 111:20]
  assign FP32Mult1_io_b = stage1Reg_2; // @[RoPEModuleFP32.scala 112:20]
  assign FP32Mult2_io_a = stage1Reg_0; // @[RoPEModuleFP32.scala 115:20]
  assign FP32Mult2_io_b = stage1Reg_3; // @[RoPEModuleFP32.scala 116:20]
  assign FP32Mult3_io_a = stage1Reg_1; // @[RoPEModuleFP32.scala 119:20]
  assign FP32Mult3_io_b = stage1Reg_3; // @[RoPEModuleFP32.scala 120:20]
  assign FP32Sub_io_a = stage2Reg_2; // @[RoPEModuleFP32.scala 132:18]
  assign FP32Sub_io_b = stage2Reg_1; // @[RoPEModuleFP32.scala 133:18]
  assign FP32add_io_a = stage2Reg_3; // @[RoPEModuleFP32.scala 136:18]
  assign FP32add_io_b = stage2Reg_0; // @[RoPEModuleFP32.scala 137:18]
  always @(posedge clock) begin
    stage1Reg_0 <= io_x_0; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_1 <= io_x_1; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_2 <= io_sin; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_3 <= io_cos; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage2Reg_0 <= FP32Mult0_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_1 <= FP32Mult1_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_2 <= FP32Mult2_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_3 <= FP32Mult3_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    if (reset) begin // @[RoPEModuleFP32.scala 97:28]
      stage3Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 97:28]
    end else begin
      stage3Reg_0 <= _WIRE_1_0; // @[RoPEModuleFP32.scala 139:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 97:28]
      stage3Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 97:28]
    end else begin
      stage3Reg_1 <= _WIRE_1_1; // @[RoPEModuleFP32.scala 139:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_0 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_0 <= io_EN; // @[RoPEModuleFP32.scala 101:14]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_1 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_1 <= enReg_0; // @[RoPEModuleFP32.scala 102:14]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_2 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_2 <= enReg_1; // @[RoPEModuleFP32.scala 103:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage1Reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage1Reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stage1Reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stage2Reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stage2Reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stage2Reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage2Reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage3Reg_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage3Reg_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  enReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  enReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  enReg_2 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP32RoPEmodule(
  input         clock,
  input         reset,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_m,
  input  [31:0] io_baseIndex,
  input  [31:0] io_TwoDivD,
  output [31:0] io_xhat_0,
  output [31:0] io_xhat_1,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  RadCacl_clock; // @[RoPEModuleFP32.scala 166:27]
  wire  RadCacl_reset; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_x_0; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_x_1; // @[RoPEModuleFP32.scala 166:27]
  wire  RadCacl_io_EN; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_m; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_baseIndex; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_TwoDivD; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_out; // @[RoPEModuleFP32.scala 166:27]
  wire  RadCacl_io_ENout; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_xFWD_0; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] RadCacl_io_xFWD_1; // @[RoPEModuleFP32.scala 166:27]
  wire [31:0] SinCosLut_io_x_0; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_x_1; // @[RoPEModuleFP32.scala 167:27]
  wire  SinCosLut_io_EN; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_angle; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_sinOut; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_cosOut; // @[RoPEModuleFP32.scala 167:27]
  wire  SinCosLut_io_ENout; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_xFWD_0; // @[RoPEModuleFP32.scala 167:27]
  wire [31:0] SinCosLut_io_xFWD_1; // @[RoPEModuleFP32.scala 167:27]
  wire  RoPEcore_clock; // @[RoPEModuleFP32.scala 168:27]
  wire  RoPEcore_reset; // @[RoPEModuleFP32.scala 168:27]
  wire  RoPEcore_io_EN; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_x_0; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_x_1; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_sin; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_cos; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_xhat_0; // @[RoPEModuleFP32.scala 168:27]
  wire [31:0] RoPEcore_io_xhat_1; // @[RoPEModuleFP32.scala 168:27]
  wire  RoPEcore_io_ENout; // @[RoPEModuleFP32.scala 168:27]
  reg [31:0] stage1Reg_0; // @[RoPEModuleFP32.scala 171:28]
  reg [31:0] stage1Reg_1; // @[RoPEModuleFP32.scala 171:28]
  reg [31:0] stage1Reg_2; // @[RoPEModuleFP32.scala 171:28]
  reg [31:0] stage1Reg_3; // @[RoPEModuleFP32.scala 171:28]
  reg [31:0] stage1Reg_4; // @[RoPEModuleFP32.scala 171:28]
  reg  stage1EN; // @[RoPEModuleFP32.scala 172:28]
  reg [31:0] stage2Reg_0; // @[RoPEModuleFP32.scala 173:28]
  reg [31:0] stage2Reg_1; // @[RoPEModuleFP32.scala 173:28]
  reg [31:0] stage2Reg_2; // @[RoPEModuleFP32.scala 173:28]
  reg  stage2EN; // @[RoPEModuleFP32.scala 174:28]
  reg [31:0] stage3Reg_0; // @[RoPEModuleFP32.scala 175:28]
  reg [31:0] stage3Reg_1; // @[RoPEModuleFP32.scala 175:28]
  reg [31:0] stage3Reg_2; // @[RoPEModuleFP32.scala 175:28]
  reg [31:0] stage3Reg_3; // @[RoPEModuleFP32.scala 175:28]
  reg  stage3EN; // @[RoPEModuleFP32.scala 176:28]
  reg [31:0] outputReg_0; // @[RoPEModuleFP32.scala 225:28]
  reg [31:0] outputReg_1; // @[RoPEModuleFP32.scala 225:28]
  reg  validReg; // @[RoPEModuleFP32.scala 226:28]
  FP32radianCaclulator RadCacl ( // @[RoPEModuleFP32.scala 166:27]
    .clock(RadCacl_clock),
    .reset(RadCacl_reset),
    .io_x_0(RadCacl_io_x_0),
    .io_x_1(RadCacl_io_x_1),
    .io_EN(RadCacl_io_EN),
    .io_m(RadCacl_io_m),
    .io_baseIndex(RadCacl_io_baseIndex),
    .io_TwoDivD(RadCacl_io_TwoDivD),
    .io_out(RadCacl_io_out),
    .io_ENout(RadCacl_io_ENout),
    .io_xFWD_0(RadCacl_io_xFWD_0),
    .io_xFWD_1(RadCacl_io_xFWD_1)
  );
  SinCosLUT SinCosLut ( // @[RoPEModuleFP32.scala 167:27]
    .io_x_0(SinCosLut_io_x_0),
    .io_x_1(SinCosLut_io_x_1),
    .io_EN(SinCosLut_io_EN),
    .io_angle(SinCosLut_io_angle),
    .io_sinOut(SinCosLut_io_sinOut),
    .io_cosOut(SinCosLut_io_cosOut),
    .io_ENout(SinCosLut_io_ENout),
    .io_xFWD_0(SinCosLut_io_xFWD_0),
    .io_xFWD_1(SinCosLut_io_xFWD_1)
  );
  FP32RoPEcore RoPEcore ( // @[RoPEModuleFP32.scala 168:27]
    .clock(RoPEcore_clock),
    .reset(RoPEcore_reset),
    .io_EN(RoPEcore_io_EN),
    .io_x_0(RoPEcore_io_x_0),
    .io_x_1(RoPEcore_io_x_1),
    .io_sin(RoPEcore_io_sin),
    .io_cos(RoPEcore_io_cos),
    .io_xhat_0(RoPEcore_io_xhat_0),
    .io_xhat_1(RoPEcore_io_xhat_1),
    .io_ENout(RoPEcore_io_ENout)
  );
  assign io_xhat_0 = outputReg_0; // @[RoPEModuleFP32.scala 228:16]
  assign io_xhat_1 = outputReg_1; // @[RoPEModuleFP32.scala 229:16]
  assign io_valid = validReg; // @[RoPEModuleFP32.scala 230:16]
  assign RadCacl_clock = clock;
  assign RadCacl_reset = reset;
  assign RadCacl_io_x_0 = stage1Reg_0; // @[RoPEModuleFP32.scala 192:29]
  assign RadCacl_io_x_1 = stage1Reg_1; // @[RoPEModuleFP32.scala 193:29]
  assign RadCacl_io_EN = stage1EN; // @[RoPEModuleFP32.scala 191:29]
  assign RadCacl_io_m = stage1Reg_2; // @[RoPEModuleFP32.scala 194:29]
  assign RadCacl_io_baseIndex = stage1Reg_3; // @[RoPEModuleFP32.scala 195:29]
  assign RadCacl_io_TwoDivD = stage1Reg_4; // @[RoPEModuleFP32.scala 196:31]
  assign SinCosLut_io_x_0 = stage2Reg_0; // @[RoPEModuleFP32.scala 207:25]
  assign SinCosLut_io_x_1 = stage2Reg_1; // @[RoPEModuleFP32.scala 208:25]
  assign SinCosLut_io_EN = stage2EN; // @[RoPEModuleFP32.scala 205:25]
  assign SinCosLut_io_angle = stage2Reg_2; // @[RoPEModuleFP32.scala 206:25]
  assign RoPEcore_clock = clock;
  assign RoPEcore_reset = reset;
  assign RoPEcore_io_EN = stage3EN; // @[RoPEModuleFP32.scala 218:25]
  assign RoPEcore_io_x_0 = stage3Reg_0; // @[RoPEModuleFP32.scala 219:25]
  assign RoPEcore_io_x_1 = stage3Reg_1; // @[RoPEModuleFP32.scala 220:25]
  assign RoPEcore_io_sin = stage3Reg_2; // @[RoPEModuleFP32.scala 221:25]
  assign RoPEcore_io_cos = stage3Reg_3; // @[RoPEModuleFP32.scala 222:25]
  always @(posedge clock) begin
    if (reset) begin // @[RoPEModuleFP32.scala 171:28]
      stage1Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 171:28]
    end else if (io_EN) begin // @[RoPEModuleFP32.scala 179:17]
      stage1Reg_0 <= io_x_0; // @[RoPEModuleFP32.scala 180:22]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 171:28]
      stage1Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 171:28]
    end else if (io_EN) begin // @[RoPEModuleFP32.scala 179:17]
      stage1Reg_1 <= io_x_1; // @[RoPEModuleFP32.scala 181:22]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 171:28]
      stage1Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 171:28]
    end else if (io_EN) begin // @[RoPEModuleFP32.scala 179:17]
      stage1Reg_2 <= io_m; // @[RoPEModuleFP32.scala 182:22]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 171:28]
      stage1Reg_3 <= 32'h0; // @[RoPEModuleFP32.scala 171:28]
    end else if (io_EN) begin // @[RoPEModuleFP32.scala 179:17]
      stage1Reg_3 <= io_baseIndex; // @[RoPEModuleFP32.scala 183:22]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 171:28]
      stage1Reg_4 <= 32'h0; // @[RoPEModuleFP32.scala 171:28]
    end else if (io_EN) begin // @[RoPEModuleFP32.scala 179:17]
      stage1Reg_4 <= io_TwoDivD; // @[RoPEModuleFP32.scala 184:22]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 172:28]
      stage1EN <= 1'h0; // @[RoPEModuleFP32.scala 172:28]
    end else begin
      stage1EN <= io_EN;
    end
    if (reset) begin // @[RoPEModuleFP32.scala 173:28]
      stage2Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 173:28]
    end else begin
      stage2Reg_0 <= RadCacl_io_xFWD_0; // @[RoPEModuleFP32.scala 199:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 173:28]
      stage2Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 173:28]
    end else begin
      stage2Reg_1 <= RadCacl_io_xFWD_1; // @[RoPEModuleFP32.scala 200:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 173:28]
      stage2Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 173:28]
    end else begin
      stage2Reg_2 <= RadCacl_io_out; // @[RoPEModuleFP32.scala 201:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 174:28]
      stage2EN <= 1'h0; // @[RoPEModuleFP32.scala 174:28]
    end else begin
      stage2EN <= RadCacl_io_ENout; // @[RoPEModuleFP32.scala 202:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 175:28]
      stage3Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 175:28]
    end else begin
      stage3Reg_0 <= SinCosLut_io_xFWD_0; // @[RoPEModuleFP32.scala 211:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 175:28]
      stage3Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 175:28]
    end else begin
      stage3Reg_1 <= SinCosLut_io_xFWD_1; // @[RoPEModuleFP32.scala 212:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 175:28]
      stage3Reg_2 <= 32'h0; // @[RoPEModuleFP32.scala 175:28]
    end else begin
      stage3Reg_2 <= SinCosLut_io_sinOut; // @[RoPEModuleFP32.scala 213:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 175:28]
      stage3Reg_3 <= 32'h0; // @[RoPEModuleFP32.scala 175:28]
    end else begin
      stage3Reg_3 <= SinCosLut_io_cosOut; // @[RoPEModuleFP32.scala 214:18]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 176:28]
      stage3EN <= 1'h0; // @[RoPEModuleFP32.scala 176:28]
    end else begin
      stage3EN <= SinCosLut_io_ENout; // @[RoPEModuleFP32.scala 215:18]
    end
    outputReg_0 <= RoPEcore_io_xhat_0; // @[RoPEModuleFP32.scala 225:{36,36}]
    outputReg_1 <= RoPEcore_io_xhat_1; // @[RoPEModuleFP32.scala 225:{36,36}]
    validReg <= RoPEcore_io_ENout; // @[RoPEModuleFP32.scala 226:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage1Reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage1Reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stage1Reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stage1Reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stage1EN = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stage2Reg_0 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage2Reg_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage2Reg_2 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage2EN = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  stage3Reg_0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stage3Reg_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stage3Reg_2 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  stage3Reg_3 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stage3EN = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  outputReg_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  outputReg_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  validReg = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
