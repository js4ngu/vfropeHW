module FP32radianCaclulatorV2(
  input         clock,
  input         reset,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_m,
  input  [31:0] io_baseIndex,
  input  [31:0] io_ResMode,
  output [31:0] io_out,
  output        io_ENout,
  output [31:0] io_xFWD_0,
  output [31:0] io_xFWD_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] _stage1Reg_T = {{1'd0}, io_baseIndex}; // @[RoPEModuleFP32v2.scala 19:73]
  wire [63:0] _stage1Reg_T_2 = io_m * _stage1Reg_T[31:0]; // @[RoPEModuleFP32v2.scala 19:57]
  wire [43:0] _stage1Reg_T_4 = io_ResMode * _stage1Reg_T_2[11:0]; // @[RoPEModuleFP32v2.scala 19:49]
  reg [31:0] stage1Reg_0; // @[RoPEModuleFP32v2.scala 18:28]
  reg [31:0] stage1Reg_1; // @[RoPEModuleFP32v2.scala 18:28]
  reg [31:0] stage1Reg_2; // @[RoPEModuleFP32v2.scala 18:28]
  reg  enReg_0; // @[RoPEModuleFP32v2.scala 21:28]
  assign io_out = enReg_0 ? stage1Reg_2 : 32'h0; // @[RoPEModuleFP32v2.scala 30:22]
  assign io_ENout = enReg_0; // @[RoPEModuleFP32v2.scala 31:16]
  assign io_xFWD_0 = enReg_0 ? stage1Reg_0 : 32'h0; // @[RoPEModuleFP32v2.scala 28:22]
  assign io_xFWD_1 = enReg_0 ? stage1Reg_1 : 32'h0; // @[RoPEModuleFP32v2.scala 29:22]
  always @(posedge clock) begin
    stage1Reg_0 <= io_x_0; // @[RoPEModuleFP32v2.scala 18:{36,36}]
    stage1Reg_1 <= io_x_1; // @[RoPEModuleFP32v2.scala 18:{36,36}]
    stage1Reg_2 <= {{20'd0}, _stage1Reg_T_4[11:0]}; // @[RoPEModuleFP32v2.scala 18:{36,36}]
    if (reset) begin // @[RoPEModuleFP32v2.scala 21:28]
      enReg_0 <= 1'h0; // @[RoPEModuleFP32v2.scala 21:28]
    end else begin
      enReg_0 <= io_EN; // @[RoPEModuleFP32v2.scala 24:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage1Reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage1Reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  enReg_0 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module decoder(
  input  [31:0] io_cosIndex1,
  input  [31:0] io_sinIndex1,
  output [31:0] io_cosIndex2,
  output [31:0] io_sinIndex2,
  output        io_cosSign,
  output        io_sinSign
);
  wire [31:0] _cosIndexWire_T_1 = 32'h800 - io_cosIndex1; // @[sincosLUT2.scala 91:30]
  wire  _T_2 = io_cosIndex1 <= 32'hc00; // @[sincosLUT2.scala 93:29]
  wire [31:0] _cosIndexWire_T_3 = io_cosIndex1 - 32'h800; // @[sincosLUT2.scala 94:38]
  wire [31:0] _cosIndexWire_T_5 = 32'h1000 - io_cosIndex1; // @[sincosLUT2.scala 97:36]
  wire [31:0] _GEN_0 = io_cosIndex1 <= 32'hc00 ? _cosIndexWire_T_3 : _cosIndexWire_T_5; // @[sincosLUT2.scala 93:48 94:22 97:22]
  wire [31:0] _GEN_2 = io_cosIndex1 <= 32'h800 ? _cosIndexWire_T_1 : _GEN_0; // @[sincosLUT2.scala 90:38 91:22]
  wire  _GEN_3 = io_cosIndex1 <= 32'h800 | _T_2; // @[sincosLUT2.scala 90:38 92:22]
  wire [31:0] _sinIndexWire_T_1 = 32'h800 - io_sinIndex1; // @[sincosLUT2.scala 105:30]
  wire [31:0] _sinIndexWire_T_3 = io_sinIndex1 - 32'h800; // @[sincosLUT2.scala 108:38]
  wire [31:0] _sinIndexWire_T_5 = 32'h1000 - io_sinIndex1; // @[sincosLUT2.scala 111:36]
  wire [31:0] _GEN_6 = io_sinIndex1 <= 32'hc00 ? _sinIndexWire_T_3 : _sinIndexWire_T_5; // @[sincosLUT2.scala 107:48 108:22 111:22]
  wire  _GEN_7 = io_sinIndex1 <= 32'hc00 ? 1'h0 : 1'h1; // @[sincosLUT2.scala 107:48 109:22 112:22]
  wire [31:0] _GEN_8 = io_sinIndex1 <= 32'h800 ? _sinIndexWire_T_1 : _GEN_6; // @[sincosLUT2.scala 104:38 105:22]
  wire  _GEN_9 = io_sinIndex1 <= 32'h800 ? 1'h0 : _GEN_7; // @[sincosLUT2.scala 104:38 106:22]
  assign io_cosIndex2 = io_cosIndex1 <= 32'h400 ? io_cosIndex1 : _GEN_2; // @[sincosLUT2.scala 87:36 88:22]
  assign io_sinIndex2 = io_sinIndex1 <= 32'h400 ? io_sinIndex1 : _GEN_8; // @[sincosLUT2.scala 101:36 102:22]
  assign io_cosSign = io_cosIndex1 <= 32'h400 ? 1'h0 : _GEN_3; // @[sincosLUT2.scala 87:36 89:22]
  assign io_sinSign = io_sinIndex1 <= 32'h400 | _GEN_9; // @[sincosLUT2.scala 101:36 103:22]
endmodule
module dualPortIndexCalculatorV2(
  input         clock,
  input         reset,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_angle,
  output [31:0] io_cosIndex,
  output [31:0] io_sinIndex,
  output        io_cosSign,
  output        io_sinSign,
  output        io_ENout,
  output [31:0] io_xFWD_0,
  output [31:0] io_xFWD_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] decoder_io_cosIndex1; // @[sincosLUT3.scala 36:25]
  wire [31:0] decoder_io_sinIndex1; // @[sincosLUT3.scala 36:25]
  wire [31:0] decoder_io_cosIndex2; // @[sincosLUT3.scala 36:25]
  wire [31:0] decoder_io_sinIndex2; // @[sincosLUT3.scala 36:25]
  wire  decoder_io_cosSign; // @[sincosLUT3.scala 36:25]
  wire  decoder_io_sinSign; // @[sincosLUT3.scala 36:25]
  reg [31:0] stage1Reg; // @[sincosLUT3.scala 20:33]
  reg [31:0] stage2Reg_0; // @[sincosLUT3.scala 21:33]
  reg [31:0] stage2Reg_1; // @[sincosLUT3.scala 21:33]
  reg [31:0] stage2Reg_2; // @[sincosLUT3.scala 21:33]
  reg [31:0] stage2Reg_3; // @[sincosLUT3.scala 21:33]
  reg [31:0] x0Reg_0; // @[sincosLUT3.scala 25:24]
  reg [31:0] x0Reg_1; // @[sincosLUT3.scala 25:24]
  reg [31:0] x1Reg_0; // @[sincosLUT3.scala 26:24]
  reg [31:0] x1Reg_1; // @[sincosLUT3.scala 26:24]
  reg  ENReg_0; // @[sincosLUT3.scala 27:24]
  reg  ENReg_1; // @[sincosLUT3.scala 27:24]
  wire [31:0] _decoder_io_sinIndex1_T_1 = stage1Reg + 32'h400; // @[sincosLUT3.scala 38:40]
  wire [31:0] _io_cosSign_T = ENReg_1 ? stage2Reg_2 : 32'h0; // @[sincosLUT3.scala 48:23]
  wire [31:0] _io_sinSign_T = ENReg_1 ? stage2Reg_3 : 32'h0; // @[sincosLUT3.scala 49:23]
  decoder decoder ( // @[sincosLUT3.scala 36:25]
    .io_cosIndex1(decoder_io_cosIndex1),
    .io_sinIndex1(decoder_io_sinIndex1),
    .io_cosIndex2(decoder_io_cosIndex2),
    .io_sinIndex2(decoder_io_sinIndex2),
    .io_cosSign(decoder_io_cosSign),
    .io_sinSign(decoder_io_sinSign)
  );
  assign io_cosIndex = ENReg_1 ? stage2Reg_0 : 32'h0; // @[sincosLUT3.scala 46:23]
  assign io_sinIndex = ENReg_1 ? stage2Reg_1 : 32'h0; // @[sincosLUT3.scala 47:23]
  assign io_cosSign = _io_cosSign_T[0]; // @[sincosLUT3.scala 48:17]
  assign io_sinSign = _io_sinSign_T[0]; // @[sincosLUT3.scala 49:17]
  assign io_ENout = ENReg_1; // @[sincosLUT3.scala 52:17]
  assign io_xFWD_0 = ENReg_1 ? x0Reg_1 : 32'h0; // @[sincosLUT3.scala 50:23]
  assign io_xFWD_1 = ENReg_1 ? x1Reg_1 : 32'h0; // @[sincosLUT3.scala 51:23]
  assign decoder_io_cosIndex1 = stage1Reg; // @[sincosLUT3.scala 37:26]
  assign decoder_io_sinIndex1 = {{20'd0}, _decoder_io_sinIndex1_T_1[11:0]}; // @[sincosLUT3.scala 38:26]
  always @(posedge clock) begin
    if (reset) begin // @[sincosLUT3.scala 20:33]
      stage1Reg <= 32'h0; // @[sincosLUT3.scala 20:33]
    end else begin
      stage1Reg <= io_angle; // @[sincosLUT3.scala 22:15]
    end
    if (reset) begin // @[sincosLUT3.scala 21:33]
      stage2Reg_0 <= 32'h0; // @[sincosLUT3.scala 21:33]
    end else begin
      stage2Reg_0 <= decoder_io_cosIndex2; // @[sincosLUT3.scala 40:18]
    end
    if (reset) begin // @[sincosLUT3.scala 21:33]
      stage2Reg_1 <= 32'h0; // @[sincosLUT3.scala 21:33]
    end else begin
      stage2Reg_1 <= decoder_io_sinIndex2; // @[sincosLUT3.scala 41:18]
    end
    if (reset) begin // @[sincosLUT3.scala 21:33]
      stage2Reg_2 <= 32'h0; // @[sincosLUT3.scala 21:33]
    end else begin
      stage2Reg_2 <= {{31'd0}, decoder_io_cosSign}; // @[sincosLUT3.scala 42:18]
    end
    if (reset) begin // @[sincosLUT3.scala 21:33]
      stage2Reg_3 <= 32'h0; // @[sincosLUT3.scala 21:33]
    end else begin
      stage2Reg_3 <= {{31'd0}, decoder_io_sinSign}; // @[sincosLUT3.scala 43:18]
    end
    if (reset) begin // @[sincosLUT3.scala 25:24]
      x0Reg_0 <= 32'h0; // @[sincosLUT3.scala 25:24]
    end else begin
      x0Reg_0 <= io_x_0; // @[sincosLUT3.scala 31:14]
    end
    if (reset) begin // @[sincosLUT3.scala 25:24]
      x0Reg_1 <= 32'h0; // @[sincosLUT3.scala 25:24]
    end else begin
      x0Reg_1 <= x0Reg_0; // @[sincosLUT3.scala 32:14]
    end
    if (reset) begin // @[sincosLUT3.scala 26:24]
      x1Reg_0 <= 32'h0; // @[sincosLUT3.scala 26:24]
    end else begin
      x1Reg_0 <= io_x_1; // @[sincosLUT3.scala 33:14]
    end
    if (reset) begin // @[sincosLUT3.scala 26:24]
      x1Reg_1 <= 32'h0; // @[sincosLUT3.scala 26:24]
    end else begin
      x1Reg_1 <= x1Reg_0; // @[sincosLUT3.scala 34:14]
    end
    if (reset) begin // @[sincosLUT3.scala 27:24]
      ENReg_0 <= 1'h0; // @[sincosLUT3.scala 27:24]
    end else begin
      ENReg_0 <= io_EN; // @[sincosLUT3.scala 29:14]
    end
    if (reset) begin // @[sincosLUT3.scala 27:24]
      ENReg_1 <= 1'h0; // @[sincosLUT3.scala 27:24]
    end else begin
      ENReg_1 <= ENReg_0; // @[sincosLUT3.scala 30:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage2Reg_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage2Reg_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stage2Reg_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stage2Reg_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  x0Reg_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  x0Reg_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  x1Reg_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  x1Reg_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  ENReg_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ENReg_1 = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multiPortCOSlut(
  input         clock,
  input         reset,
  input         io_EN,
  input  [31:0] io_x_0_0,
  input  [31:0] io_x_0_1,
  input  [31:0] io_x_1_0,
  input  [31:0] io_x_1_1,
  input  [31:0] io_x_2_0,
  input  [31:0] io_x_2_1,
  input  [31:0] io_x_3_0,
  input  [31:0] io_x_3_1,
  input  [31:0] io_x_4_0,
  input  [31:0] io_x_4_1,
  input  [31:0] io_x_5_0,
  input  [31:0] io_x_5_1,
  input  [31:0] io_x_6_0,
  input  [31:0] io_x_6_1,
  input  [31:0] io_x_7_0,
  input  [31:0] io_x_7_1,
  input  [31:0] io_cosIndex_0,
  input  [31:0] io_cosIndex_1,
  input  [31:0] io_cosIndex_2,
  input  [31:0] io_cosIndex_3,
  input  [31:0] io_cosIndex_4,
  input  [31:0] io_cosIndex_5,
  input  [31:0] io_cosIndex_6,
  input  [31:0] io_cosIndex_7,
  input  [31:0] io_sinIndex_0,
  input  [31:0] io_sinIndex_1,
  input  [31:0] io_sinIndex_2,
  input  [31:0] io_sinIndex_3,
  input  [31:0] io_sinIndex_4,
  input  [31:0] io_sinIndex_5,
  input  [31:0] io_sinIndex_6,
  input  [31:0] io_sinIndex_7,
  input         io_sign_0_0,
  input         io_sign_0_1,
  input         io_sign_1_0,
  input         io_sign_1_1,
  input         io_sign_2_0,
  input         io_sign_2_1,
  input         io_sign_3_0,
  input         io_sign_3_1,
  input         io_sign_4_0,
  input         io_sign_4_1,
  input         io_sign_5_0,
  input         io_sign_5_1,
  input         io_sign_6_0,
  input         io_sign_6_1,
  input         io_sign_7_0,
  input         io_sign_7_1,
  output [31:0] io_sinOut_0,
  output [31:0] io_sinOut_1,
  output [31:0] io_sinOut_2,
  output [31:0] io_sinOut_3,
  output [31:0] io_sinOut_4,
  output [31:0] io_sinOut_5,
  output [31:0] io_sinOut_6,
  output [31:0] io_sinOut_7,
  output [31:0] io_cosOut_0,
  output [31:0] io_cosOut_1,
  output [31:0] io_cosOut_2,
  output [31:0] io_cosOut_3,
  output [31:0] io_cosOut_4,
  output [31:0] io_cosOut_5,
  output [31:0] io_cosOut_6,
  output [31:0] io_cosOut_7,
  output        io_ENout,
  output [31:0] io_xFWD_0_0,
  output [31:0] io_xFWD_0_1,
  output [31:0] io_xFWD_1_0,
  output [31:0] io_xFWD_1_1,
  output [31:0] io_xFWD_2_0,
  output [31:0] io_xFWD_2_1,
  output [31:0] io_xFWD_3_0,
  output [31:0] io_xFWD_3_1,
  output [31:0] io_xFWD_4_0,
  output [31:0] io_xFWD_4_1,
  output [31:0] io_xFWD_5_0,
  output [31:0] io_xFWD_5_1,
  output [31:0] io_xFWD_6_0,
  output [31:0] io_xFWD_6_1,
  output [31:0] io_xFWD_7_0,
  output [31:0] io_xFWD_7_1,
  output        io_signFWD_0_0,
  output        io_signFWD_0_1,
  output        io_signFWD_1_0,
  output        io_signFWD_1_1,
  output        io_signFWD_2_0,
  output        io_signFWD_2_1,
  output        io_signFWD_3_0,
  output        io_signFWD_3_1,
  output        io_signFWD_4_0,
  output        io_signFWD_4_1,
  output        io_signFWD_5_0,
  output        io_signFWD_5_1,
  output        io_signFWD_6_0,
  output        io_signFWD_6_1,
  output        io_signFWD_7_0,
  output        io_signFWD_7_1
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cosLUT [0:1024]; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_0_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_0_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_0_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_0_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_0_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_0_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_1_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_1_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_1_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_1_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_1_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_1_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_2_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_2_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_2_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_2_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_2_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_2_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_3_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_3_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_3_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_3_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_3_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_3_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_4_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_4_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_4_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_4_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_4_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_4_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_5_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_5_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_5_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_5_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_5_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_5_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_6_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_6_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_6_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_6_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_6_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_6_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_cosOut_7_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_cosOut_7_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_cosOut_7_MPORT_data; // @[LUTbank2.scala 323:29]
  wire  cosLUT_io_sinOut_7_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_io_sinOut_7_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_io_sinOut_7_MPORT_data; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_2_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_2_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_2_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_2_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_3_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_3_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_3_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_3_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_4_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_4_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_4_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_4_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_5_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_5_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_5_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_5_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_6_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_6_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_6_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_6_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_7_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_7_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_7_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_7_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_8_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_8_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_8_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_8_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_9_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_9_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_9_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_9_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_10_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_10_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_10_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_10_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_11_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_11_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_11_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_11_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_12_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_12_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_12_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_12_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_13_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_13_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_13_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_13_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_14_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_14_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_14_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_14_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_15_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_15_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_15_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_15_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_16_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_16_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_16_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_16_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_17_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_17_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_17_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_17_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_18_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_18_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_18_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_18_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_19_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_19_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_19_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_19_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_20_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_20_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_20_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_20_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_21_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_21_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_21_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_21_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_22_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_22_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_22_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_22_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_23_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_23_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_23_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_23_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_24_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_24_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_24_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_24_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_25_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_25_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_25_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_25_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_26_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_26_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_26_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_26_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_27_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_27_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_27_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_27_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_28_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_28_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_28_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_28_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_29_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_29_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_29_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_29_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_30_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_30_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_30_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_30_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_31_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_31_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_31_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_31_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_32_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_32_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_32_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_32_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_33_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_33_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_33_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_33_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_34_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_34_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_34_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_34_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_35_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_35_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_35_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_35_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_36_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_36_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_36_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_36_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_37_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_37_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_37_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_37_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_38_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_38_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_38_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_38_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_39_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_39_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_39_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_39_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_40_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_40_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_40_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_40_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_41_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_41_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_41_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_41_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_42_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_42_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_42_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_42_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_43_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_43_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_43_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_43_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_44_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_44_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_44_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_44_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_45_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_45_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_45_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_45_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_46_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_46_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_46_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_46_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_47_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_47_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_47_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_47_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_48_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_48_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_48_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_48_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_49_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_49_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_49_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_49_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_50_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_50_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_50_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_50_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_51_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_51_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_51_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_51_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_52_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_52_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_52_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_52_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_53_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_53_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_53_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_53_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_54_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_54_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_54_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_54_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_55_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_55_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_55_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_55_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_56_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_56_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_56_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_56_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_57_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_57_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_57_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_57_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_58_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_58_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_58_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_58_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_59_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_59_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_59_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_59_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_60_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_60_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_60_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_60_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_61_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_61_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_61_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_61_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_62_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_62_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_62_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_62_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_63_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_63_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_63_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_63_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_64_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_64_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_64_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_64_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_65_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_65_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_65_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_65_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_66_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_66_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_66_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_66_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_67_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_67_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_67_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_67_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_68_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_68_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_68_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_68_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_69_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_69_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_69_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_69_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_70_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_70_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_70_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_70_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_71_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_71_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_71_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_71_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_72_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_72_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_72_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_72_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_73_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_73_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_73_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_73_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_74_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_74_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_74_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_74_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_75_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_75_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_75_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_75_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_76_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_76_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_76_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_76_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_77_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_77_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_77_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_77_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_78_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_78_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_78_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_78_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_79_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_79_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_79_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_79_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_80_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_80_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_80_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_80_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_81_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_81_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_81_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_81_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_82_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_82_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_82_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_82_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_83_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_83_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_83_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_83_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_84_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_84_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_84_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_84_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_85_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_85_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_85_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_85_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_86_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_86_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_86_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_86_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_87_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_87_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_87_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_87_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_88_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_88_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_88_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_88_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_89_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_89_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_89_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_89_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_90_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_90_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_90_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_90_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_91_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_91_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_91_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_91_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_92_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_92_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_92_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_92_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_93_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_93_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_93_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_93_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_94_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_94_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_94_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_94_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_95_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_95_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_95_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_95_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_96_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_96_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_96_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_96_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_97_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_97_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_97_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_97_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_98_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_98_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_98_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_98_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_99_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_99_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_99_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_99_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_100_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_100_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_100_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_100_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_101_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_101_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_101_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_101_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_102_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_102_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_102_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_102_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_103_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_103_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_103_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_103_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_104_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_104_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_104_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_104_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_105_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_105_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_105_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_105_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_106_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_106_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_106_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_106_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_107_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_107_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_107_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_107_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_108_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_108_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_108_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_108_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_109_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_109_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_109_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_109_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_110_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_110_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_110_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_110_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_111_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_111_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_111_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_111_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_112_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_112_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_112_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_112_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_113_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_113_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_113_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_113_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_114_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_114_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_114_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_114_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_115_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_115_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_115_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_115_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_116_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_116_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_116_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_116_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_117_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_117_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_117_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_117_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_118_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_118_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_118_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_118_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_119_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_119_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_119_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_119_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_120_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_120_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_120_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_120_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_121_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_121_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_121_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_121_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_122_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_122_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_122_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_122_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_123_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_123_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_123_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_123_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_124_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_124_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_124_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_124_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_125_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_125_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_125_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_125_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_126_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_126_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_126_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_126_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_127_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_127_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_127_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_127_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_128_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_128_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_128_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_128_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_129_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_129_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_129_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_129_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_130_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_130_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_130_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_130_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_131_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_131_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_131_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_131_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_132_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_132_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_132_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_132_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_133_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_133_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_133_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_133_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_134_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_134_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_134_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_134_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_135_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_135_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_135_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_135_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_136_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_136_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_136_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_136_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_137_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_137_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_137_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_137_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_138_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_138_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_138_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_138_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_139_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_139_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_139_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_139_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_140_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_140_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_140_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_140_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_141_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_141_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_141_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_141_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_142_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_142_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_142_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_142_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_143_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_143_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_143_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_143_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_144_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_144_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_144_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_144_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_145_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_145_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_145_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_145_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_146_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_146_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_146_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_146_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_147_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_147_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_147_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_147_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_148_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_148_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_148_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_148_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_149_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_149_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_149_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_149_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_150_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_150_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_150_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_150_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_151_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_151_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_151_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_151_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_152_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_152_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_152_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_152_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_153_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_153_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_153_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_153_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_154_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_154_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_154_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_154_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_155_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_155_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_155_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_155_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_156_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_156_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_156_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_156_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_157_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_157_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_157_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_157_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_158_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_158_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_158_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_158_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_159_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_159_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_159_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_159_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_160_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_160_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_160_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_160_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_161_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_161_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_161_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_161_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_162_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_162_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_162_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_162_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_163_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_163_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_163_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_163_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_164_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_164_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_164_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_164_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_165_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_165_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_165_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_165_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_166_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_166_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_166_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_166_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_167_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_167_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_167_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_167_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_168_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_168_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_168_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_168_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_169_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_169_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_169_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_169_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_170_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_170_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_170_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_170_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_171_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_171_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_171_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_171_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_172_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_172_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_172_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_172_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_173_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_173_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_173_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_173_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_174_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_174_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_174_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_174_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_175_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_175_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_175_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_175_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_176_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_176_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_176_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_176_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_177_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_177_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_177_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_177_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_178_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_178_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_178_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_178_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_179_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_179_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_179_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_179_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_180_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_180_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_180_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_180_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_181_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_181_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_181_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_181_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_182_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_182_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_182_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_182_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_183_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_183_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_183_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_183_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_184_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_184_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_184_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_184_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_185_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_185_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_185_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_185_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_186_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_186_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_186_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_186_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_187_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_187_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_187_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_187_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_188_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_188_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_188_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_188_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_189_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_189_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_189_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_189_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_190_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_190_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_190_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_190_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_191_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_191_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_191_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_191_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_192_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_192_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_192_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_192_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_193_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_193_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_193_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_193_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_194_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_194_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_194_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_194_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_195_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_195_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_195_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_195_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_196_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_196_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_196_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_196_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_197_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_197_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_197_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_197_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_198_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_198_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_198_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_198_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_199_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_199_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_199_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_199_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_200_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_200_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_200_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_200_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_201_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_201_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_201_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_201_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_202_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_202_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_202_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_202_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_203_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_203_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_203_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_203_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_204_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_204_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_204_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_204_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_205_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_205_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_205_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_205_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_206_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_206_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_206_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_206_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_207_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_207_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_207_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_207_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_208_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_208_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_208_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_208_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_209_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_209_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_209_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_209_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_210_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_210_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_210_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_210_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_211_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_211_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_211_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_211_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_212_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_212_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_212_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_212_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_213_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_213_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_213_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_213_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_214_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_214_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_214_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_214_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_215_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_215_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_215_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_215_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_216_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_216_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_216_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_216_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_217_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_217_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_217_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_217_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_218_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_218_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_218_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_218_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_219_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_219_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_219_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_219_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_220_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_220_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_220_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_220_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_221_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_221_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_221_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_221_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_222_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_222_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_222_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_222_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_223_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_223_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_223_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_223_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_224_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_224_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_224_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_224_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_225_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_225_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_225_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_225_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_226_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_226_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_226_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_226_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_227_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_227_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_227_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_227_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_228_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_228_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_228_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_228_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_229_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_229_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_229_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_229_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_230_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_230_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_230_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_230_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_231_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_231_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_231_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_231_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_232_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_232_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_232_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_232_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_233_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_233_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_233_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_233_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_234_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_234_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_234_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_234_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_235_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_235_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_235_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_235_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_236_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_236_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_236_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_236_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_237_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_237_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_237_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_237_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_238_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_238_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_238_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_238_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_239_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_239_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_239_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_239_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_240_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_240_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_240_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_240_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_241_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_241_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_241_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_241_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_242_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_242_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_242_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_242_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_243_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_243_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_243_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_243_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_244_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_244_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_244_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_244_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_245_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_245_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_245_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_245_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_246_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_246_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_246_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_246_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_247_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_247_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_247_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_247_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_248_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_248_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_248_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_248_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_249_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_249_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_249_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_249_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_250_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_250_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_250_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_250_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_251_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_251_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_251_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_251_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_252_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_252_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_252_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_252_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_253_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_253_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_253_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_253_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_254_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_254_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_254_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_254_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_255_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_255_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_255_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_255_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_256_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_256_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_256_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_256_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_257_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_257_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_257_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_257_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_258_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_258_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_258_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_258_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_259_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_259_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_259_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_259_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_260_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_260_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_260_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_260_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_261_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_261_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_261_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_261_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_262_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_262_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_262_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_262_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_263_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_263_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_263_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_263_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_264_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_264_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_264_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_264_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_265_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_265_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_265_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_265_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_266_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_266_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_266_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_266_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_267_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_267_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_267_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_267_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_268_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_268_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_268_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_268_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_269_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_269_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_269_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_269_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_270_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_270_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_270_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_270_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_271_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_271_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_271_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_271_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_272_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_272_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_272_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_272_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_273_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_273_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_273_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_273_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_274_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_274_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_274_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_274_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_275_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_275_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_275_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_275_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_276_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_276_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_276_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_276_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_277_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_277_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_277_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_277_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_278_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_278_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_278_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_278_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_279_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_279_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_279_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_279_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_280_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_280_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_280_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_280_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_281_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_281_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_281_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_281_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_282_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_282_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_282_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_282_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_283_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_283_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_283_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_283_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_284_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_284_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_284_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_284_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_285_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_285_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_285_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_285_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_286_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_286_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_286_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_286_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_287_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_287_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_287_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_287_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_288_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_288_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_288_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_288_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_289_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_289_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_289_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_289_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_290_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_290_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_290_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_290_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_291_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_291_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_291_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_291_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_292_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_292_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_292_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_292_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_293_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_293_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_293_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_293_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_294_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_294_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_294_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_294_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_295_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_295_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_295_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_295_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_296_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_296_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_296_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_296_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_297_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_297_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_297_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_297_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_298_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_298_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_298_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_298_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_299_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_299_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_299_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_299_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_300_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_300_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_300_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_300_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_301_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_301_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_301_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_301_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_302_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_302_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_302_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_302_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_303_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_303_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_303_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_303_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_304_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_304_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_304_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_304_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_305_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_305_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_305_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_305_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_306_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_306_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_306_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_306_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_307_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_307_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_307_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_307_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_308_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_308_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_308_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_308_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_309_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_309_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_309_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_309_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_310_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_310_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_310_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_310_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_311_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_311_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_311_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_311_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_312_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_312_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_312_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_312_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_313_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_313_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_313_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_313_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_314_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_314_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_314_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_314_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_315_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_315_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_315_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_315_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_316_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_316_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_316_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_316_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_317_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_317_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_317_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_317_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_318_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_318_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_318_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_318_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_319_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_319_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_319_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_319_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_320_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_320_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_320_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_320_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_321_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_321_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_321_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_321_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_322_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_322_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_322_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_322_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_323_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_323_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_323_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_323_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_324_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_324_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_324_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_324_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_325_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_325_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_325_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_325_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_326_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_326_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_326_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_326_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_327_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_327_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_327_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_327_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_328_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_328_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_328_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_328_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_329_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_329_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_329_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_329_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_330_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_330_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_330_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_330_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_331_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_331_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_331_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_331_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_332_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_332_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_332_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_332_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_333_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_333_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_333_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_333_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_334_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_334_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_334_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_334_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_335_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_335_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_335_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_335_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_336_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_336_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_336_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_336_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_337_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_337_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_337_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_337_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_338_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_338_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_338_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_338_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_339_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_339_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_339_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_339_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_340_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_340_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_340_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_340_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_341_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_341_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_341_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_341_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_342_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_342_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_342_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_342_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_343_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_343_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_343_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_343_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_344_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_344_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_344_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_344_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_345_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_345_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_345_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_345_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_346_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_346_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_346_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_346_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_347_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_347_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_347_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_347_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_348_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_348_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_348_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_348_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_349_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_349_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_349_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_349_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_350_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_350_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_350_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_350_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_351_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_351_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_351_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_351_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_352_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_352_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_352_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_352_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_353_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_353_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_353_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_353_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_354_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_354_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_354_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_354_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_355_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_355_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_355_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_355_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_356_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_356_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_356_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_356_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_357_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_357_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_357_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_357_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_358_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_358_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_358_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_358_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_359_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_359_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_359_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_359_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_360_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_360_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_360_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_360_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_361_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_361_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_361_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_361_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_362_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_362_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_362_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_362_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_363_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_363_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_363_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_363_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_364_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_364_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_364_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_364_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_365_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_365_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_365_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_365_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_366_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_366_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_366_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_366_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_367_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_367_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_367_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_367_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_368_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_368_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_368_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_368_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_369_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_369_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_369_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_369_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_370_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_370_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_370_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_370_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_371_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_371_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_371_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_371_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_372_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_372_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_372_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_372_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_373_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_373_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_373_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_373_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_374_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_374_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_374_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_374_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_375_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_375_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_375_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_375_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_376_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_376_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_376_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_376_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_377_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_377_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_377_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_377_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_378_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_378_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_378_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_378_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_379_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_379_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_379_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_379_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_380_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_380_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_380_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_380_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_381_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_381_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_381_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_381_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_382_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_382_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_382_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_382_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_383_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_383_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_383_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_383_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_384_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_384_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_384_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_384_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_385_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_385_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_385_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_385_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_386_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_386_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_386_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_386_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_387_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_387_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_387_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_387_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_388_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_388_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_388_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_388_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_389_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_389_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_389_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_389_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_390_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_390_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_390_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_390_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_391_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_391_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_391_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_391_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_392_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_392_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_392_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_392_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_393_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_393_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_393_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_393_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_394_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_394_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_394_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_394_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_395_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_395_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_395_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_395_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_396_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_396_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_396_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_396_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_397_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_397_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_397_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_397_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_398_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_398_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_398_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_398_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_399_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_399_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_399_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_399_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_400_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_400_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_400_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_400_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_401_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_401_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_401_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_401_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_402_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_402_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_402_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_402_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_403_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_403_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_403_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_403_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_404_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_404_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_404_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_404_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_405_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_405_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_405_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_405_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_406_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_406_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_406_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_406_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_407_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_407_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_407_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_407_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_408_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_408_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_408_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_408_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_409_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_409_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_409_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_409_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_410_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_410_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_410_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_410_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_411_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_411_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_411_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_411_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_412_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_412_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_412_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_412_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_413_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_413_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_413_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_413_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_414_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_414_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_414_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_414_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_415_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_415_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_415_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_415_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_416_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_416_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_416_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_416_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_417_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_417_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_417_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_417_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_418_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_418_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_418_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_418_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_419_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_419_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_419_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_419_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_420_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_420_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_420_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_420_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_421_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_421_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_421_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_421_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_422_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_422_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_422_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_422_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_423_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_423_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_423_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_423_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_424_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_424_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_424_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_424_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_425_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_425_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_425_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_425_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_426_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_426_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_426_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_426_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_427_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_427_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_427_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_427_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_428_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_428_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_428_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_428_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_429_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_429_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_429_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_429_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_430_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_430_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_430_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_430_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_431_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_431_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_431_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_431_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_432_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_432_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_432_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_432_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_433_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_433_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_433_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_433_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_434_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_434_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_434_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_434_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_435_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_435_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_435_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_435_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_436_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_436_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_436_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_436_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_437_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_437_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_437_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_437_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_438_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_438_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_438_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_438_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_439_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_439_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_439_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_439_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_440_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_440_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_440_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_440_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_441_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_441_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_441_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_441_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_442_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_442_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_442_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_442_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_443_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_443_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_443_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_443_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_444_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_444_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_444_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_444_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_445_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_445_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_445_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_445_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_446_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_446_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_446_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_446_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_447_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_447_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_447_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_447_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_448_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_448_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_448_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_448_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_449_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_449_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_449_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_449_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_450_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_450_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_450_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_450_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_451_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_451_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_451_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_451_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_452_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_452_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_452_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_452_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_453_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_453_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_453_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_453_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_454_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_454_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_454_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_454_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_455_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_455_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_455_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_455_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_456_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_456_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_456_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_456_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_457_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_457_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_457_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_457_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_458_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_458_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_458_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_458_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_459_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_459_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_459_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_459_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_460_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_460_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_460_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_460_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_461_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_461_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_461_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_461_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_462_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_462_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_462_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_462_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_463_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_463_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_463_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_463_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_464_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_464_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_464_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_464_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_465_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_465_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_465_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_465_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_466_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_466_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_466_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_466_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_467_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_467_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_467_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_467_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_468_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_468_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_468_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_468_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_469_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_469_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_469_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_469_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_470_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_470_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_470_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_470_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_471_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_471_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_471_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_471_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_472_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_472_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_472_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_472_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_473_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_473_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_473_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_473_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_474_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_474_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_474_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_474_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_475_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_475_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_475_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_475_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_476_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_476_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_476_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_476_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_477_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_477_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_477_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_477_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_478_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_478_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_478_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_478_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_479_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_479_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_479_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_479_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_480_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_480_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_480_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_480_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_481_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_481_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_481_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_481_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_482_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_482_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_482_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_482_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_483_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_483_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_483_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_483_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_484_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_484_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_484_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_484_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_485_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_485_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_485_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_485_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_486_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_486_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_486_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_486_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_487_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_487_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_487_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_487_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_488_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_488_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_488_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_488_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_489_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_489_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_489_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_489_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_490_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_490_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_490_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_490_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_491_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_491_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_491_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_491_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_492_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_492_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_492_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_492_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_493_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_493_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_493_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_493_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_494_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_494_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_494_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_494_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_495_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_495_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_495_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_495_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_496_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_496_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_496_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_496_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_497_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_497_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_497_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_497_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_498_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_498_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_498_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_498_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_499_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_499_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_499_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_499_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_500_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_500_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_500_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_500_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_501_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_501_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_501_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_501_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_502_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_502_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_502_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_502_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_503_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_503_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_503_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_503_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_504_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_504_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_504_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_504_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_505_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_505_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_505_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_505_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_506_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_506_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_506_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_506_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_507_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_507_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_507_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_507_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_508_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_508_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_508_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_508_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_509_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_509_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_509_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_509_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_510_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_510_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_510_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_510_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_511_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_511_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_511_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_511_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_512_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_512_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_512_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_512_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_513_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_513_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_513_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_513_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_514_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_514_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_514_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_514_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_515_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_515_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_515_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_515_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_516_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_516_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_516_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_516_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_517_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_517_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_517_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_517_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_518_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_518_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_518_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_518_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_519_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_519_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_519_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_519_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_520_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_520_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_520_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_520_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_521_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_521_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_521_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_521_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_522_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_522_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_522_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_522_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_523_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_523_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_523_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_523_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_524_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_524_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_524_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_524_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_525_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_525_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_525_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_525_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_526_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_526_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_526_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_526_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_527_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_527_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_527_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_527_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_528_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_528_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_528_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_528_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_529_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_529_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_529_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_529_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_530_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_530_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_530_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_530_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_531_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_531_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_531_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_531_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_532_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_532_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_532_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_532_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_533_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_533_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_533_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_533_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_534_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_534_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_534_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_534_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_535_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_535_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_535_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_535_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_536_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_536_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_536_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_536_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_537_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_537_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_537_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_537_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_538_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_538_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_538_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_538_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_539_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_539_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_539_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_539_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_540_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_540_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_540_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_540_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_541_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_541_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_541_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_541_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_542_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_542_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_542_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_542_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_543_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_543_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_543_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_543_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_544_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_544_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_544_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_544_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_545_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_545_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_545_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_545_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_546_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_546_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_546_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_546_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_547_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_547_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_547_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_547_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_548_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_548_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_548_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_548_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_549_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_549_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_549_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_549_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_550_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_550_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_550_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_550_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_551_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_551_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_551_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_551_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_552_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_552_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_552_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_552_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_553_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_553_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_553_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_553_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_554_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_554_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_554_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_554_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_555_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_555_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_555_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_555_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_556_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_556_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_556_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_556_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_557_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_557_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_557_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_557_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_558_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_558_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_558_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_558_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_559_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_559_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_559_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_559_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_560_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_560_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_560_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_560_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_561_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_561_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_561_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_561_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_562_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_562_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_562_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_562_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_563_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_563_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_563_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_563_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_564_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_564_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_564_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_564_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_565_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_565_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_565_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_565_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_566_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_566_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_566_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_566_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_567_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_567_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_567_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_567_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_568_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_568_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_568_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_568_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_569_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_569_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_569_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_569_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_570_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_570_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_570_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_570_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_571_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_571_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_571_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_571_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_572_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_572_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_572_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_572_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_573_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_573_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_573_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_573_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_574_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_574_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_574_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_574_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_575_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_575_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_575_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_575_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_576_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_576_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_576_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_576_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_577_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_577_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_577_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_577_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_578_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_578_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_578_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_578_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_579_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_579_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_579_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_579_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_580_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_580_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_580_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_580_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_581_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_581_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_581_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_581_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_582_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_582_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_582_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_582_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_583_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_583_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_583_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_583_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_584_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_584_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_584_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_584_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_585_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_585_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_585_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_585_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_586_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_586_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_586_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_586_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_587_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_587_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_587_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_587_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_588_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_588_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_588_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_588_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_589_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_589_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_589_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_589_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_590_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_590_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_590_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_590_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_591_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_591_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_591_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_591_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_592_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_592_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_592_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_592_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_593_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_593_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_593_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_593_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_594_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_594_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_594_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_594_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_595_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_595_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_595_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_595_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_596_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_596_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_596_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_596_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_597_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_597_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_597_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_597_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_598_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_598_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_598_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_598_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_599_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_599_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_599_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_599_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_600_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_600_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_600_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_600_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_601_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_601_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_601_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_601_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_602_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_602_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_602_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_602_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_603_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_603_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_603_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_603_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_604_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_604_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_604_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_604_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_605_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_605_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_605_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_605_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_606_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_606_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_606_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_606_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_607_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_607_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_607_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_607_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_608_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_608_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_608_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_608_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_609_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_609_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_609_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_609_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_610_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_610_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_610_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_610_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_611_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_611_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_611_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_611_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_612_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_612_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_612_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_612_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_613_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_613_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_613_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_613_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_614_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_614_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_614_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_614_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_615_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_615_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_615_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_615_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_616_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_616_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_616_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_616_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_617_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_617_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_617_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_617_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_618_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_618_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_618_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_618_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_619_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_619_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_619_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_619_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_620_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_620_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_620_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_620_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_621_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_621_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_621_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_621_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_622_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_622_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_622_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_622_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_623_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_623_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_623_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_623_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_624_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_624_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_624_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_624_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_625_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_625_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_625_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_625_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_626_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_626_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_626_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_626_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_627_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_627_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_627_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_627_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_628_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_628_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_628_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_628_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_629_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_629_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_629_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_629_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_630_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_630_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_630_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_630_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_631_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_631_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_631_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_631_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_632_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_632_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_632_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_632_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_633_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_633_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_633_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_633_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_634_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_634_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_634_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_634_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_635_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_635_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_635_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_635_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_636_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_636_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_636_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_636_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_637_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_637_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_637_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_637_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_638_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_638_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_638_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_638_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_639_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_639_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_639_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_639_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_640_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_640_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_640_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_640_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_641_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_641_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_641_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_641_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_642_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_642_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_642_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_642_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_643_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_643_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_643_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_643_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_644_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_644_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_644_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_644_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_645_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_645_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_645_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_645_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_646_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_646_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_646_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_646_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_647_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_647_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_647_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_647_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_648_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_648_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_648_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_648_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_649_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_649_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_649_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_649_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_650_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_650_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_650_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_650_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_651_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_651_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_651_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_651_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_652_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_652_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_652_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_652_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_653_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_653_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_653_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_653_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_654_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_654_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_654_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_654_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_655_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_655_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_655_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_655_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_656_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_656_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_656_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_656_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_657_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_657_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_657_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_657_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_658_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_658_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_658_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_658_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_659_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_659_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_659_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_659_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_660_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_660_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_660_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_660_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_661_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_661_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_661_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_661_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_662_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_662_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_662_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_662_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_663_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_663_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_663_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_663_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_664_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_664_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_664_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_664_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_665_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_665_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_665_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_665_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_666_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_666_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_666_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_666_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_667_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_667_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_667_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_667_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_668_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_668_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_668_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_668_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_669_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_669_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_669_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_669_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_670_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_670_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_670_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_670_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_671_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_671_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_671_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_671_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_672_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_672_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_672_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_672_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_673_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_673_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_673_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_673_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_674_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_674_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_674_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_674_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_675_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_675_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_675_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_675_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_676_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_676_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_676_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_676_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_677_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_677_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_677_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_677_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_678_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_678_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_678_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_678_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_679_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_679_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_679_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_679_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_680_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_680_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_680_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_680_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_681_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_681_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_681_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_681_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_682_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_682_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_682_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_682_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_683_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_683_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_683_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_683_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_684_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_684_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_684_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_684_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_685_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_685_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_685_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_685_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_686_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_686_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_686_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_686_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_687_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_687_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_687_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_687_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_688_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_688_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_688_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_688_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_689_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_689_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_689_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_689_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_690_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_690_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_690_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_690_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_691_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_691_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_691_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_691_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_692_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_692_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_692_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_692_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_693_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_693_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_693_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_693_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_694_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_694_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_694_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_694_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_695_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_695_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_695_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_695_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_696_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_696_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_696_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_696_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_697_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_697_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_697_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_697_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_698_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_698_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_698_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_698_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_699_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_699_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_699_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_699_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_700_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_700_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_700_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_700_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_701_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_701_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_701_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_701_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_702_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_702_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_702_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_702_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_703_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_703_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_703_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_703_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_704_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_704_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_704_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_704_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_705_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_705_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_705_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_705_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_706_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_706_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_706_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_706_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_707_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_707_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_707_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_707_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_708_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_708_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_708_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_708_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_709_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_709_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_709_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_709_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_710_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_710_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_710_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_710_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_711_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_711_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_711_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_711_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_712_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_712_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_712_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_712_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_713_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_713_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_713_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_713_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_714_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_714_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_714_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_714_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_715_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_715_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_715_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_715_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_716_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_716_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_716_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_716_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_717_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_717_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_717_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_717_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_718_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_718_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_718_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_718_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_719_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_719_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_719_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_719_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_720_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_720_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_720_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_720_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_721_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_721_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_721_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_721_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_722_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_722_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_722_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_722_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_723_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_723_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_723_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_723_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_724_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_724_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_724_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_724_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_725_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_725_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_725_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_725_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_726_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_726_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_726_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_726_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_727_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_727_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_727_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_727_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_728_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_728_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_728_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_728_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_729_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_729_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_729_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_729_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_730_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_730_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_730_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_730_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_731_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_731_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_731_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_731_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_732_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_732_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_732_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_732_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_733_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_733_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_733_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_733_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_734_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_734_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_734_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_734_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_735_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_735_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_735_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_735_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_736_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_736_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_736_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_736_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_737_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_737_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_737_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_737_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_738_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_738_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_738_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_738_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_739_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_739_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_739_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_739_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_740_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_740_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_740_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_740_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_741_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_741_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_741_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_741_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_742_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_742_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_742_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_742_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_743_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_743_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_743_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_743_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_744_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_744_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_744_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_744_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_745_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_745_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_745_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_745_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_746_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_746_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_746_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_746_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_747_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_747_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_747_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_747_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_748_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_748_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_748_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_748_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_749_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_749_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_749_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_749_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_750_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_750_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_750_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_750_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_751_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_751_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_751_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_751_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_752_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_752_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_752_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_752_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_753_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_753_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_753_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_753_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_754_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_754_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_754_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_754_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_755_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_755_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_755_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_755_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_756_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_756_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_756_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_756_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_757_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_757_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_757_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_757_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_758_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_758_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_758_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_758_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_759_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_759_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_759_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_759_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_760_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_760_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_760_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_760_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_761_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_761_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_761_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_761_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_762_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_762_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_762_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_762_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_763_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_763_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_763_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_763_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_764_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_764_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_764_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_764_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_765_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_765_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_765_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_765_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_766_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_766_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_766_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_766_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_767_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_767_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_767_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_767_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_768_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_768_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_768_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_768_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_769_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_769_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_769_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_769_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_770_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_770_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_770_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_770_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_771_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_771_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_771_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_771_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_772_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_772_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_772_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_772_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_773_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_773_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_773_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_773_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_774_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_774_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_774_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_774_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_775_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_775_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_775_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_775_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_776_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_776_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_776_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_776_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_777_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_777_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_777_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_777_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_778_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_778_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_778_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_778_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_779_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_779_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_779_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_779_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_780_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_780_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_780_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_780_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_781_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_781_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_781_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_781_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_782_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_782_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_782_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_782_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_783_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_783_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_783_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_783_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_784_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_784_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_784_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_784_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_785_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_785_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_785_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_785_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_786_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_786_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_786_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_786_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_787_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_787_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_787_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_787_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_788_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_788_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_788_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_788_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_789_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_789_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_789_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_789_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_790_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_790_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_790_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_790_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_791_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_791_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_791_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_791_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_792_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_792_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_792_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_792_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_793_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_793_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_793_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_793_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_794_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_794_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_794_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_794_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_795_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_795_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_795_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_795_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_796_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_796_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_796_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_796_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_797_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_797_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_797_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_797_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_798_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_798_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_798_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_798_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_799_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_799_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_799_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_799_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_800_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_800_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_800_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_800_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_801_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_801_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_801_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_801_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_802_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_802_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_802_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_802_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_803_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_803_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_803_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_803_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_804_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_804_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_804_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_804_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_805_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_805_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_805_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_805_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_806_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_806_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_806_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_806_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_807_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_807_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_807_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_807_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_808_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_808_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_808_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_808_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_809_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_809_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_809_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_809_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_810_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_810_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_810_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_810_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_811_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_811_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_811_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_811_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_812_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_812_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_812_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_812_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_813_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_813_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_813_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_813_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_814_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_814_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_814_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_814_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_815_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_815_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_815_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_815_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_816_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_816_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_816_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_816_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_817_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_817_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_817_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_817_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_818_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_818_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_818_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_818_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_819_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_819_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_819_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_819_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_820_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_820_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_820_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_820_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_821_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_821_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_821_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_821_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_822_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_822_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_822_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_822_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_823_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_823_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_823_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_823_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_824_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_824_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_824_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_824_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_825_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_825_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_825_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_825_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_826_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_826_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_826_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_826_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_827_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_827_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_827_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_827_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_828_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_828_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_828_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_828_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_829_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_829_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_829_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_829_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_830_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_830_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_830_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_830_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_831_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_831_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_831_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_831_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_832_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_832_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_832_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_832_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_833_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_833_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_833_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_833_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_834_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_834_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_834_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_834_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_835_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_835_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_835_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_835_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_836_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_836_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_836_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_836_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_837_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_837_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_837_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_837_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_838_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_838_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_838_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_838_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_839_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_839_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_839_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_839_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_840_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_840_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_840_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_840_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_841_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_841_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_841_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_841_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_842_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_842_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_842_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_842_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_843_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_843_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_843_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_843_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_844_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_844_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_844_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_844_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_845_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_845_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_845_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_845_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_846_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_846_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_846_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_846_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_847_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_847_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_847_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_847_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_848_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_848_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_848_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_848_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_849_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_849_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_849_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_849_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_850_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_850_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_850_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_850_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_851_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_851_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_851_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_851_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_852_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_852_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_852_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_852_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_853_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_853_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_853_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_853_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_854_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_854_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_854_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_854_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_855_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_855_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_855_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_855_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_856_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_856_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_856_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_856_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_857_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_857_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_857_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_857_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_858_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_858_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_858_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_858_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_859_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_859_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_859_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_859_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_860_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_860_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_860_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_860_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_861_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_861_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_861_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_861_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_862_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_862_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_862_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_862_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_863_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_863_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_863_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_863_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_864_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_864_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_864_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_864_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_865_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_865_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_865_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_865_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_866_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_866_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_866_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_866_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_867_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_867_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_867_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_867_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_868_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_868_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_868_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_868_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_869_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_869_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_869_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_869_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_870_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_870_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_870_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_870_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_871_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_871_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_871_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_871_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_872_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_872_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_872_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_872_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_873_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_873_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_873_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_873_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_874_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_874_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_874_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_874_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_875_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_875_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_875_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_875_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_876_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_876_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_876_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_876_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_877_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_877_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_877_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_877_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_878_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_878_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_878_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_878_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_879_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_879_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_879_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_879_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_880_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_880_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_880_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_880_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_881_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_881_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_881_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_881_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_882_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_882_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_882_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_882_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_883_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_883_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_883_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_883_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_884_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_884_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_884_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_884_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_885_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_885_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_885_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_885_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_886_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_886_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_886_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_886_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_887_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_887_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_887_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_887_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_888_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_888_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_888_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_888_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_889_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_889_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_889_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_889_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_890_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_890_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_890_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_890_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_891_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_891_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_891_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_891_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_892_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_892_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_892_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_892_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_893_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_893_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_893_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_893_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_894_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_894_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_894_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_894_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_895_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_895_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_895_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_895_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_896_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_896_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_896_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_896_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_897_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_897_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_897_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_897_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_898_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_898_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_898_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_898_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_899_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_899_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_899_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_899_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_900_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_900_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_900_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_900_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_901_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_901_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_901_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_901_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_902_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_902_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_902_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_902_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_903_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_903_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_903_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_903_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_904_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_904_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_904_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_904_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_905_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_905_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_905_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_905_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_906_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_906_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_906_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_906_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_907_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_907_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_907_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_907_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_908_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_908_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_908_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_908_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_909_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_909_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_909_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_909_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_910_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_910_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_910_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_910_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_911_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_911_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_911_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_911_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_912_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_912_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_912_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_912_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_913_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_913_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_913_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_913_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_914_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_914_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_914_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_914_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_915_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_915_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_915_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_915_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_916_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_916_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_916_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_916_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_917_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_917_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_917_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_917_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_918_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_918_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_918_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_918_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_919_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_919_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_919_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_919_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_920_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_920_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_920_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_920_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_921_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_921_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_921_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_921_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_922_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_922_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_922_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_922_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_923_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_923_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_923_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_923_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_924_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_924_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_924_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_924_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_925_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_925_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_925_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_925_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_926_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_926_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_926_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_926_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_927_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_927_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_927_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_927_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_928_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_928_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_928_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_928_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_929_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_929_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_929_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_929_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_930_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_930_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_930_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_930_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_931_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_931_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_931_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_931_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_932_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_932_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_932_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_932_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_933_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_933_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_933_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_933_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_934_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_934_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_934_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_934_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_935_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_935_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_935_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_935_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_936_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_936_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_936_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_936_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_937_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_937_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_937_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_937_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_938_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_938_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_938_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_938_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_939_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_939_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_939_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_939_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_940_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_940_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_940_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_940_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_941_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_941_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_941_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_941_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_942_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_942_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_942_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_942_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_943_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_943_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_943_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_943_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_944_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_944_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_944_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_944_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_945_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_945_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_945_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_945_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_946_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_946_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_946_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_946_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_947_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_947_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_947_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_947_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_948_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_948_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_948_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_948_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_949_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_949_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_949_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_949_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_950_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_950_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_950_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_950_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_951_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_951_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_951_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_951_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_952_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_952_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_952_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_952_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_953_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_953_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_953_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_953_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_954_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_954_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_954_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_954_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_955_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_955_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_955_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_955_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_956_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_956_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_956_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_956_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_957_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_957_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_957_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_957_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_958_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_958_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_958_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_958_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_959_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_959_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_959_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_959_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_960_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_960_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_960_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_960_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_961_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_961_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_961_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_961_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_962_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_962_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_962_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_962_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_963_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_963_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_963_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_963_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_964_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_964_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_964_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_964_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_965_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_965_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_965_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_965_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_966_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_966_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_966_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_966_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_967_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_967_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_967_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_967_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_968_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_968_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_968_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_968_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_969_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_969_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_969_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_969_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_970_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_970_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_970_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_970_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_971_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_971_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_971_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_971_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_972_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_972_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_972_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_972_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_973_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_973_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_973_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_973_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_974_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_974_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_974_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_974_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_975_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_975_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_975_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_975_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_976_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_976_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_976_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_976_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_977_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_977_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_977_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_977_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_978_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_978_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_978_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_978_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_979_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_979_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_979_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_979_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_980_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_980_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_980_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_980_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_981_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_981_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_981_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_981_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_982_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_982_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_982_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_982_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_983_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_983_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_983_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_983_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_984_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_984_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_984_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_984_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_985_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_985_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_985_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_985_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_986_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_986_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_986_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_986_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_987_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_987_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_987_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_987_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_988_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_988_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_988_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_988_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_989_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_989_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_989_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_989_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_990_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_990_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_990_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_990_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_991_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_991_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_991_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_991_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_992_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_992_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_992_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_992_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_993_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_993_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_993_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_993_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_994_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_994_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_994_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_994_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_995_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_995_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_995_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_995_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_996_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_996_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_996_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_996_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_997_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_997_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_997_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_997_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_998_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_998_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_998_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_998_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_999_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_999_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_999_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_999_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1000_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1000_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1000_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1000_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1001_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1001_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1001_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1001_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1002_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1002_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1002_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1002_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1003_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1003_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1003_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1003_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1004_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1004_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1004_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1004_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1005_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1005_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1005_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1005_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1006_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1006_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1006_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1006_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1007_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1007_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1007_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1007_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1008_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1008_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1008_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1008_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1009_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1009_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1009_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1009_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1010_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1010_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1010_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1010_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1011_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1011_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1011_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1011_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1012_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1012_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1012_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1012_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1013_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1013_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1013_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1013_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1014_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1014_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1014_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1014_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1015_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1015_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1015_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1015_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1016_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1016_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1016_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1016_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1017_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1017_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1017_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1017_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1018_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1018_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1018_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1018_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1019_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1019_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1019_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1019_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1020_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1020_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1020_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1020_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1021_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1021_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1021_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1021_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1022_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1022_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1022_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1022_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1023_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1023_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1023_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1023_en; // @[LUTbank2.scala 323:29]
  wire [31:0] cosLUT_MPORT_1024_data; // @[LUTbank2.scala 323:29]
  wire [10:0] cosLUT_MPORT_1024_addr; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1024_mask; // @[LUTbank2.scala 323:29]
  wire  cosLUT_MPORT_1024_en; // @[LUTbank2.scala 323:29]
  reg  cosLUT_io_cosOut_0_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_0_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_0_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_0_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_1_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_1_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_1_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_1_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_2_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_2_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_2_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_2_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_3_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_3_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_3_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_3_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_4_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_4_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_4_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_4_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_5_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_5_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_5_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_5_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_6_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_6_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_6_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_6_MPORT_addr_pipe_0;
  reg  cosLUT_io_cosOut_7_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_cosOut_7_MPORT_addr_pipe_0;
  reg  cosLUT_io_sinOut_7_MPORT_en_pipe_0;
  reg [10:0] cosLUT_io_sinOut_7_MPORT_addr_pipe_0;
  reg  ENReg; // @[LUTbank2.scala 331:29]
  reg [31:0] xFWDReg_0_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_0_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_1_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_1_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_2_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_2_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_3_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_3_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_4_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_4_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_5_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_5_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_6_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_6_1; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_7_0; // @[LUTbank2.scala 332:29]
  reg [31:0] xFWDReg_7_1; // @[LUTbank2.scala 332:29]
  reg  signReg_0_0; // @[LUTbank2.scala 333:29]
  reg  signReg_0_1; // @[LUTbank2.scala 333:29]
  reg  signReg_1_0; // @[LUTbank2.scala 333:29]
  reg  signReg_1_1; // @[LUTbank2.scala 333:29]
  reg  signReg_2_0; // @[LUTbank2.scala 333:29]
  reg  signReg_2_1; // @[LUTbank2.scala 333:29]
  reg  signReg_3_0; // @[LUTbank2.scala 333:29]
  reg  signReg_3_1; // @[LUTbank2.scala 333:29]
  reg  signReg_4_0; // @[LUTbank2.scala 333:29]
  reg  signReg_4_1; // @[LUTbank2.scala 333:29]
  reg  signReg_5_0; // @[LUTbank2.scala 333:29]
  reg  signReg_5_1; // @[LUTbank2.scala 333:29]
  reg  signReg_6_0; // @[LUTbank2.scala 333:29]
  reg  signReg_6_1; // @[LUTbank2.scala 333:29]
  reg  signReg_7_0; // @[LUTbank2.scala 333:29]
  reg  signReg_7_1; // @[LUTbank2.scala 333:29]
  assign cosLUT_io_cosOut_0_MPORT_en = cosLUT_io_cosOut_0_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_0_MPORT_addr = cosLUT_io_cosOut_0_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_0_MPORT_data = cosLUT[cosLUT_io_cosOut_0_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_0_MPORT_data = cosLUT_io_cosOut_0_MPORT_addr >= 11'h401 ? _RAND_1[31:0] :
    cosLUT[cosLUT_io_cosOut_0_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_0_MPORT_en = cosLUT_io_sinOut_0_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_0_MPORT_addr = cosLUT_io_sinOut_0_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_0_MPORT_data = cosLUT[cosLUT_io_sinOut_0_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_0_MPORT_data = cosLUT_io_sinOut_0_MPORT_addr >= 11'h401 ? _RAND_2[31:0] :
    cosLUT[cosLUT_io_sinOut_0_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_1_MPORT_en = cosLUT_io_cosOut_1_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_1_MPORT_addr = cosLUT_io_cosOut_1_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_1_MPORT_data = cosLUT[cosLUT_io_cosOut_1_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_1_MPORT_data = cosLUT_io_cosOut_1_MPORT_addr >= 11'h401 ? _RAND_3[31:0] :
    cosLUT[cosLUT_io_cosOut_1_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_1_MPORT_en = cosLUT_io_sinOut_1_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_1_MPORT_addr = cosLUT_io_sinOut_1_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_1_MPORT_data = cosLUT[cosLUT_io_sinOut_1_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_1_MPORT_data = cosLUT_io_sinOut_1_MPORT_addr >= 11'h401 ? _RAND_4[31:0] :
    cosLUT[cosLUT_io_sinOut_1_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_2_MPORT_en = cosLUT_io_cosOut_2_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_2_MPORT_addr = cosLUT_io_cosOut_2_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_2_MPORT_data = cosLUT[cosLUT_io_cosOut_2_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_2_MPORT_data = cosLUT_io_cosOut_2_MPORT_addr >= 11'h401 ? _RAND_5[31:0] :
    cosLUT[cosLUT_io_cosOut_2_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_2_MPORT_en = cosLUT_io_sinOut_2_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_2_MPORT_addr = cosLUT_io_sinOut_2_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_2_MPORT_data = cosLUT[cosLUT_io_sinOut_2_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_2_MPORT_data = cosLUT_io_sinOut_2_MPORT_addr >= 11'h401 ? _RAND_6[31:0] :
    cosLUT[cosLUT_io_sinOut_2_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_3_MPORT_en = cosLUT_io_cosOut_3_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_3_MPORT_addr = cosLUT_io_cosOut_3_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_3_MPORT_data = cosLUT[cosLUT_io_cosOut_3_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_3_MPORT_data = cosLUT_io_cosOut_3_MPORT_addr >= 11'h401 ? _RAND_7[31:0] :
    cosLUT[cosLUT_io_cosOut_3_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_3_MPORT_en = cosLUT_io_sinOut_3_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_3_MPORT_addr = cosLUT_io_sinOut_3_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_3_MPORT_data = cosLUT[cosLUT_io_sinOut_3_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_3_MPORT_data = cosLUT_io_sinOut_3_MPORT_addr >= 11'h401 ? _RAND_8[31:0] :
    cosLUT[cosLUT_io_sinOut_3_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_4_MPORT_en = cosLUT_io_cosOut_4_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_4_MPORT_addr = cosLUT_io_cosOut_4_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_4_MPORT_data = cosLUT[cosLUT_io_cosOut_4_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_4_MPORT_data = cosLUT_io_cosOut_4_MPORT_addr >= 11'h401 ? _RAND_9[31:0] :
    cosLUT[cosLUT_io_cosOut_4_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_4_MPORT_en = cosLUT_io_sinOut_4_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_4_MPORT_addr = cosLUT_io_sinOut_4_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_4_MPORT_data = cosLUT[cosLUT_io_sinOut_4_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_4_MPORT_data = cosLUT_io_sinOut_4_MPORT_addr >= 11'h401 ? _RAND_10[31:0] :
    cosLUT[cosLUT_io_sinOut_4_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_5_MPORT_en = cosLUT_io_cosOut_5_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_5_MPORT_addr = cosLUT_io_cosOut_5_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_5_MPORT_data = cosLUT[cosLUT_io_cosOut_5_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_5_MPORT_data = cosLUT_io_cosOut_5_MPORT_addr >= 11'h401 ? _RAND_11[31:0] :
    cosLUT[cosLUT_io_cosOut_5_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_5_MPORT_en = cosLUT_io_sinOut_5_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_5_MPORT_addr = cosLUT_io_sinOut_5_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_5_MPORT_data = cosLUT[cosLUT_io_sinOut_5_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_5_MPORT_data = cosLUT_io_sinOut_5_MPORT_addr >= 11'h401 ? _RAND_12[31:0] :
    cosLUT[cosLUT_io_sinOut_5_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_6_MPORT_en = cosLUT_io_cosOut_6_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_6_MPORT_addr = cosLUT_io_cosOut_6_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_6_MPORT_data = cosLUT[cosLUT_io_cosOut_6_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_6_MPORT_data = cosLUT_io_cosOut_6_MPORT_addr >= 11'h401 ? _RAND_13[31:0] :
    cosLUT[cosLUT_io_cosOut_6_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_6_MPORT_en = cosLUT_io_sinOut_6_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_6_MPORT_addr = cosLUT_io_sinOut_6_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_6_MPORT_data = cosLUT[cosLUT_io_sinOut_6_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_6_MPORT_data = cosLUT_io_sinOut_6_MPORT_addr >= 11'h401 ? _RAND_14[31:0] :
    cosLUT[cosLUT_io_sinOut_6_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_7_MPORT_en = cosLUT_io_cosOut_7_MPORT_en_pipe_0;
  assign cosLUT_io_cosOut_7_MPORT_addr = cosLUT_io_cosOut_7_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_cosOut_7_MPORT_data = cosLUT[cosLUT_io_cosOut_7_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_cosOut_7_MPORT_data = cosLUT_io_cosOut_7_MPORT_addr >= 11'h401 ? _RAND_15[31:0] :
    cosLUT[cosLUT_io_cosOut_7_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_7_MPORT_en = cosLUT_io_sinOut_7_MPORT_en_pipe_0;
  assign cosLUT_io_sinOut_7_MPORT_addr = cosLUT_io_sinOut_7_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_io_sinOut_7_MPORT_data = cosLUT[cosLUT_io_sinOut_7_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `else
  assign cosLUT_io_sinOut_7_MPORT_data = cosLUT_io_sinOut_7_MPORT_addr >= 11'h401 ? _RAND_16[31:0] :
    cosLUT[cosLUT_io_sinOut_7_MPORT_addr]; // @[LUTbank2.scala 323:29]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosLUT_MPORT_data = 32'h3f800000;
  assign cosLUT_MPORT_addr = 11'h0;
  assign cosLUT_MPORT_mask = 1'h1;
  assign cosLUT_MPORT_en = reset;
  assign cosLUT_MPORT_1_data = 32'h3f7fffec;
  assign cosLUT_MPORT_1_addr = 11'h1;
  assign cosLUT_MPORT_1_mask = 1'h1;
  assign cosLUT_MPORT_1_en = reset;
  assign cosLUT_MPORT_2_data = 32'h3f7fffb1;
  assign cosLUT_MPORT_2_addr = 11'h2;
  assign cosLUT_MPORT_2_mask = 1'h1;
  assign cosLUT_MPORT_2_en = reset;
  assign cosLUT_MPORT_3_data = 32'h3f7fff4e;
  assign cosLUT_MPORT_3_addr = 11'h3;
  assign cosLUT_MPORT_3_mask = 1'h1;
  assign cosLUT_MPORT_3_en = reset;
  assign cosLUT_MPORT_4_data = 32'h3f7ffec4;
  assign cosLUT_MPORT_4_addr = 11'h4;
  assign cosLUT_MPORT_4_mask = 1'h1;
  assign cosLUT_MPORT_4_en = reset;
  assign cosLUT_MPORT_5_data = 32'h3f7ffe12;
  assign cosLUT_MPORT_5_addr = 11'h5;
  assign cosLUT_MPORT_5_mask = 1'h1;
  assign cosLUT_MPORT_5_en = reset;
  assign cosLUT_MPORT_6_data = 32'h3f7ffd39;
  assign cosLUT_MPORT_6_addr = 11'h6;
  assign cosLUT_MPORT_6_mask = 1'h1;
  assign cosLUT_MPORT_6_en = reset;
  assign cosLUT_MPORT_7_data = 32'h3f7ffc38;
  assign cosLUT_MPORT_7_addr = 11'h7;
  assign cosLUT_MPORT_7_mask = 1'h1;
  assign cosLUT_MPORT_7_en = reset;
  assign cosLUT_MPORT_8_data = 32'h3f7ffb10;
  assign cosLUT_MPORT_8_addr = 11'h8;
  assign cosLUT_MPORT_8_mask = 1'h1;
  assign cosLUT_MPORT_8_en = reset;
  assign cosLUT_MPORT_9_data = 32'h3f7ff9c0;
  assign cosLUT_MPORT_9_addr = 11'h9;
  assign cosLUT_MPORT_9_mask = 1'h1;
  assign cosLUT_MPORT_9_en = reset;
  assign cosLUT_MPORT_10_data = 32'h3f7ff849;
  assign cosLUT_MPORT_10_addr = 11'ha;
  assign cosLUT_MPORT_10_mask = 1'h1;
  assign cosLUT_MPORT_10_en = reset;
  assign cosLUT_MPORT_11_data = 32'h3f7ff6aa;
  assign cosLUT_MPORT_11_addr = 11'hb;
  assign cosLUT_MPORT_11_mask = 1'h1;
  assign cosLUT_MPORT_11_en = reset;
  assign cosLUT_MPORT_12_data = 32'h3f7ff4e4;
  assign cosLUT_MPORT_12_addr = 11'hc;
  assign cosLUT_MPORT_12_mask = 1'h1;
  assign cosLUT_MPORT_12_en = reset;
  assign cosLUT_MPORT_13_data = 32'h3f7ff2f7;
  assign cosLUT_MPORT_13_addr = 11'hd;
  assign cosLUT_MPORT_13_mask = 1'h1;
  assign cosLUT_MPORT_13_en = reset;
  assign cosLUT_MPORT_14_data = 32'h3f7ff0e1;
  assign cosLUT_MPORT_14_addr = 11'he;
  assign cosLUT_MPORT_14_mask = 1'h1;
  assign cosLUT_MPORT_14_en = reset;
  assign cosLUT_MPORT_15_data = 32'h3f7feea5;
  assign cosLUT_MPORT_15_addr = 11'hf;
  assign cosLUT_MPORT_15_mask = 1'h1;
  assign cosLUT_MPORT_15_en = reset;
  assign cosLUT_MPORT_16_data = 32'h3f7fec41;
  assign cosLUT_MPORT_16_addr = 11'h10;
  assign cosLUT_MPORT_16_mask = 1'h1;
  assign cosLUT_MPORT_16_en = reset;
  assign cosLUT_MPORT_17_data = 32'h3f7fe9b5;
  assign cosLUT_MPORT_17_addr = 11'h11;
  assign cosLUT_MPORT_17_mask = 1'h1;
  assign cosLUT_MPORT_17_en = reset;
  assign cosLUT_MPORT_18_data = 32'h3f7fe702;
  assign cosLUT_MPORT_18_addr = 11'h12;
  assign cosLUT_MPORT_18_mask = 1'h1;
  assign cosLUT_MPORT_18_en = reset;
  assign cosLUT_MPORT_19_data = 32'h3f7fe427;
  assign cosLUT_MPORT_19_addr = 11'h13;
  assign cosLUT_MPORT_19_mask = 1'h1;
  assign cosLUT_MPORT_19_en = reset;
  assign cosLUT_MPORT_20_data = 32'h3f7fe125;
  assign cosLUT_MPORT_20_addr = 11'h14;
  assign cosLUT_MPORT_20_mask = 1'h1;
  assign cosLUT_MPORT_20_en = reset;
  assign cosLUT_MPORT_21_data = 32'h3f7fddfc;
  assign cosLUT_MPORT_21_addr = 11'h15;
  assign cosLUT_MPORT_21_mask = 1'h1;
  assign cosLUT_MPORT_21_en = reset;
  assign cosLUT_MPORT_22_data = 32'h3f7fdaaa;
  assign cosLUT_MPORT_22_addr = 11'h16;
  assign cosLUT_MPORT_22_mask = 1'h1;
  assign cosLUT_MPORT_22_en = reset;
  assign cosLUT_MPORT_23_data = 32'h3f7fd732;
  assign cosLUT_MPORT_23_addr = 11'h17;
  assign cosLUT_MPORT_23_mask = 1'h1;
  assign cosLUT_MPORT_23_en = reset;
  assign cosLUT_MPORT_24_data = 32'h3f7fd392;
  assign cosLUT_MPORT_24_addr = 11'h18;
  assign cosLUT_MPORT_24_mask = 1'h1;
  assign cosLUT_MPORT_24_en = reset;
  assign cosLUT_MPORT_25_data = 32'h3f7fcfca;
  assign cosLUT_MPORT_25_addr = 11'h19;
  assign cosLUT_MPORT_25_mask = 1'h1;
  assign cosLUT_MPORT_25_en = reset;
  assign cosLUT_MPORT_26_data = 32'h3f7fcbdc;
  assign cosLUT_MPORT_26_addr = 11'h1a;
  assign cosLUT_MPORT_26_mask = 1'h1;
  assign cosLUT_MPORT_26_en = reset;
  assign cosLUT_MPORT_27_data = 32'h3f7fc7c5;
  assign cosLUT_MPORT_27_addr = 11'h1b;
  assign cosLUT_MPORT_27_mask = 1'h1;
  assign cosLUT_MPORT_27_en = reset;
  assign cosLUT_MPORT_28_data = 32'h3f7fc387;
  assign cosLUT_MPORT_28_addr = 11'h1c;
  assign cosLUT_MPORT_28_mask = 1'h1;
  assign cosLUT_MPORT_28_en = reset;
  assign cosLUT_MPORT_29_data = 32'h3f7fbf22;
  assign cosLUT_MPORT_29_addr = 11'h1d;
  assign cosLUT_MPORT_29_mask = 1'h1;
  assign cosLUT_MPORT_29_en = reset;
  assign cosLUT_MPORT_30_data = 32'h3f7fba95;
  assign cosLUT_MPORT_30_addr = 11'h1e;
  assign cosLUT_MPORT_30_mask = 1'h1;
  assign cosLUT_MPORT_30_en = reset;
  assign cosLUT_MPORT_31_data = 32'h3f7fb5e1;
  assign cosLUT_MPORT_31_addr = 11'h1f;
  assign cosLUT_MPORT_31_mask = 1'h1;
  assign cosLUT_MPORT_31_en = reset;
  assign cosLUT_MPORT_32_data = 32'h3f7fb105;
  assign cosLUT_MPORT_32_addr = 11'h20;
  assign cosLUT_MPORT_32_mask = 1'h1;
  assign cosLUT_MPORT_32_en = reset;
  assign cosLUT_MPORT_33_data = 32'h3f7fac02;
  assign cosLUT_MPORT_33_addr = 11'h21;
  assign cosLUT_MPORT_33_mask = 1'h1;
  assign cosLUT_MPORT_33_en = reset;
  assign cosLUT_MPORT_34_data = 32'h3f7fa6d8;
  assign cosLUT_MPORT_34_addr = 11'h22;
  assign cosLUT_MPORT_34_mask = 1'h1;
  assign cosLUT_MPORT_34_en = reset;
  assign cosLUT_MPORT_35_data = 32'h3f7fa185;
  assign cosLUT_MPORT_35_addr = 11'h23;
  assign cosLUT_MPORT_35_mask = 1'h1;
  assign cosLUT_MPORT_35_en = reset;
  assign cosLUT_MPORT_36_data = 32'h3f7f9c0c;
  assign cosLUT_MPORT_36_addr = 11'h24;
  assign cosLUT_MPORT_36_mask = 1'h1;
  assign cosLUT_MPORT_36_en = reset;
  assign cosLUT_MPORT_37_data = 32'h3f7f966b;
  assign cosLUT_MPORT_37_addr = 11'h25;
  assign cosLUT_MPORT_37_mask = 1'h1;
  assign cosLUT_MPORT_37_en = reset;
  assign cosLUT_MPORT_38_data = 32'h3f7f90a3;
  assign cosLUT_MPORT_38_addr = 11'h26;
  assign cosLUT_MPORT_38_mask = 1'h1;
  assign cosLUT_MPORT_38_en = reset;
  assign cosLUT_MPORT_39_data = 32'h3f7f8ab3;
  assign cosLUT_MPORT_39_addr = 11'h27;
  assign cosLUT_MPORT_39_mask = 1'h1;
  assign cosLUT_MPORT_39_en = reset;
  assign cosLUT_MPORT_40_data = 32'h3f7f849c;
  assign cosLUT_MPORT_40_addr = 11'h28;
  assign cosLUT_MPORT_40_mask = 1'h1;
  assign cosLUT_MPORT_40_en = reset;
  assign cosLUT_MPORT_41_data = 32'h3f7f7e5d;
  assign cosLUT_MPORT_41_addr = 11'h29;
  assign cosLUT_MPORT_41_mask = 1'h1;
  assign cosLUT_MPORT_41_en = reset;
  assign cosLUT_MPORT_42_data = 32'h3f7f77f7;
  assign cosLUT_MPORT_42_addr = 11'h2a;
  assign cosLUT_MPORT_42_mask = 1'h1;
  assign cosLUT_MPORT_42_en = reset;
  assign cosLUT_MPORT_43_data = 32'h3f7f716a;
  assign cosLUT_MPORT_43_addr = 11'h2b;
  assign cosLUT_MPORT_43_mask = 1'h1;
  assign cosLUT_MPORT_43_en = reset;
  assign cosLUT_MPORT_44_data = 32'h3f7f6ab5;
  assign cosLUT_MPORT_44_addr = 11'h2c;
  assign cosLUT_MPORT_44_mask = 1'h1;
  assign cosLUT_MPORT_44_en = reset;
  assign cosLUT_MPORT_45_data = 32'h3f7f63d8;
  assign cosLUT_MPORT_45_addr = 11'h2d;
  assign cosLUT_MPORT_45_mask = 1'h1;
  assign cosLUT_MPORT_45_en = reset;
  assign cosLUT_MPORT_46_data = 32'h3f7f5cd5;
  assign cosLUT_MPORT_46_addr = 11'h2e;
  assign cosLUT_MPORT_46_mask = 1'h1;
  assign cosLUT_MPORT_46_en = reset;
  assign cosLUT_MPORT_47_data = 32'h3f7f55aa;
  assign cosLUT_MPORT_47_addr = 11'h2f;
  assign cosLUT_MPORT_47_mask = 1'h1;
  assign cosLUT_MPORT_47_en = reset;
  assign cosLUT_MPORT_48_data = 32'h3f7f4e57;
  assign cosLUT_MPORT_48_addr = 11'h30;
  assign cosLUT_MPORT_48_mask = 1'h1;
  assign cosLUT_MPORT_48_en = reset;
  assign cosLUT_MPORT_49_data = 32'h3f7f46dd;
  assign cosLUT_MPORT_49_addr = 11'h31;
  assign cosLUT_MPORT_49_mask = 1'h1;
  assign cosLUT_MPORT_49_en = reset;
  assign cosLUT_MPORT_50_data = 32'h3f7f3f3c;
  assign cosLUT_MPORT_50_addr = 11'h32;
  assign cosLUT_MPORT_50_mask = 1'h1;
  assign cosLUT_MPORT_50_en = reset;
  assign cosLUT_MPORT_51_data = 32'h3f7f3773;
  assign cosLUT_MPORT_51_addr = 11'h33;
  assign cosLUT_MPORT_51_mask = 1'h1;
  assign cosLUT_MPORT_51_en = reset;
  assign cosLUT_MPORT_52_data = 32'h3f7f2f83;
  assign cosLUT_MPORT_52_addr = 11'h34;
  assign cosLUT_MPORT_52_mask = 1'h1;
  assign cosLUT_MPORT_52_en = reset;
  assign cosLUT_MPORT_53_data = 32'h3f7f276c;
  assign cosLUT_MPORT_53_addr = 11'h35;
  assign cosLUT_MPORT_53_mask = 1'h1;
  assign cosLUT_MPORT_53_en = reset;
  assign cosLUT_MPORT_54_data = 32'h3f7f1f2d;
  assign cosLUT_MPORT_54_addr = 11'h36;
  assign cosLUT_MPORT_54_mask = 1'h1;
  assign cosLUT_MPORT_54_en = reset;
  assign cosLUT_MPORT_55_data = 32'h3f7f16c7;
  assign cosLUT_MPORT_55_addr = 11'h37;
  assign cosLUT_MPORT_55_mask = 1'h1;
  assign cosLUT_MPORT_55_en = reset;
  assign cosLUT_MPORT_56_data = 32'h3f7f0e3a;
  assign cosLUT_MPORT_56_addr = 11'h38;
  assign cosLUT_MPORT_56_mask = 1'h1;
  assign cosLUT_MPORT_56_en = reset;
  assign cosLUT_MPORT_57_data = 32'h3f7f0585;
  assign cosLUT_MPORT_57_addr = 11'h39;
  assign cosLUT_MPORT_57_mask = 1'h1;
  assign cosLUT_MPORT_57_en = reset;
  assign cosLUT_MPORT_58_data = 32'h3f7efca9;
  assign cosLUT_MPORT_58_addr = 11'h3a;
  assign cosLUT_MPORT_58_mask = 1'h1;
  assign cosLUT_MPORT_58_en = reset;
  assign cosLUT_MPORT_59_data = 32'h3f7ef3a5;
  assign cosLUT_MPORT_59_addr = 11'h3b;
  assign cosLUT_MPORT_59_mask = 1'h1;
  assign cosLUT_MPORT_59_en = reset;
  assign cosLUT_MPORT_60_data = 32'h3f7eea7a;
  assign cosLUT_MPORT_60_addr = 11'h3c;
  assign cosLUT_MPORT_60_mask = 1'h1;
  assign cosLUT_MPORT_60_en = reset;
  assign cosLUT_MPORT_61_data = 32'h3f7ee128;
  assign cosLUT_MPORT_61_addr = 11'h3d;
  assign cosLUT_MPORT_61_mask = 1'h1;
  assign cosLUT_MPORT_61_en = reset;
  assign cosLUT_MPORT_62_data = 32'h3f7ed7af;
  assign cosLUT_MPORT_62_addr = 11'h3e;
  assign cosLUT_MPORT_62_mask = 1'h1;
  assign cosLUT_MPORT_62_en = reset;
  assign cosLUT_MPORT_63_data = 32'h3f7ece0e;
  assign cosLUT_MPORT_63_addr = 11'h3f;
  assign cosLUT_MPORT_63_mask = 1'h1;
  assign cosLUT_MPORT_63_en = reset;
  assign cosLUT_MPORT_64_data = 32'h3f7ec446;
  assign cosLUT_MPORT_64_addr = 11'h40;
  assign cosLUT_MPORT_64_mask = 1'h1;
  assign cosLUT_MPORT_64_en = reset;
  assign cosLUT_MPORT_65_data = 32'h3f7eba56;
  assign cosLUT_MPORT_65_addr = 11'h41;
  assign cosLUT_MPORT_65_mask = 1'h1;
  assign cosLUT_MPORT_65_en = reset;
  assign cosLUT_MPORT_66_data = 32'h3f7eb03f;
  assign cosLUT_MPORT_66_addr = 11'h42;
  assign cosLUT_MPORT_66_mask = 1'h1;
  assign cosLUT_MPORT_66_en = reset;
  assign cosLUT_MPORT_67_data = 32'h3f7ea601;
  assign cosLUT_MPORT_67_addr = 11'h43;
  assign cosLUT_MPORT_67_mask = 1'h1;
  assign cosLUT_MPORT_67_en = reset;
  assign cosLUT_MPORT_68_data = 32'h3f7e9b9c;
  assign cosLUT_MPORT_68_addr = 11'h44;
  assign cosLUT_MPORT_68_mask = 1'h1;
  assign cosLUT_MPORT_68_en = reset;
  assign cosLUT_MPORT_69_data = 32'h3f7e9110;
  assign cosLUT_MPORT_69_addr = 11'h45;
  assign cosLUT_MPORT_69_mask = 1'h1;
  assign cosLUT_MPORT_69_en = reset;
  assign cosLUT_MPORT_70_data = 32'h3f7e865c;
  assign cosLUT_MPORT_70_addr = 11'h46;
  assign cosLUT_MPORT_70_mask = 1'h1;
  assign cosLUT_MPORT_70_en = reset;
  assign cosLUT_MPORT_71_data = 32'h3f7e7b80;
  assign cosLUT_MPORT_71_addr = 11'h47;
  assign cosLUT_MPORT_71_mask = 1'h1;
  assign cosLUT_MPORT_71_en = reset;
  assign cosLUT_MPORT_72_data = 32'h3f7e707e;
  assign cosLUT_MPORT_72_addr = 11'h48;
  assign cosLUT_MPORT_72_mask = 1'h1;
  assign cosLUT_MPORT_72_en = reset;
  assign cosLUT_MPORT_73_data = 32'h3f7e6554;
  assign cosLUT_MPORT_73_addr = 11'h49;
  assign cosLUT_MPORT_73_mask = 1'h1;
  assign cosLUT_MPORT_73_en = reset;
  assign cosLUT_MPORT_74_data = 32'h3f7e5a03;
  assign cosLUT_MPORT_74_addr = 11'h4a;
  assign cosLUT_MPORT_74_mask = 1'h1;
  assign cosLUT_MPORT_74_en = reset;
  assign cosLUT_MPORT_75_data = 32'h3f7e4e8b;
  assign cosLUT_MPORT_75_addr = 11'h4b;
  assign cosLUT_MPORT_75_mask = 1'h1;
  assign cosLUT_MPORT_75_en = reset;
  assign cosLUT_MPORT_76_data = 32'h3f7e42ec;
  assign cosLUT_MPORT_76_addr = 11'h4c;
  assign cosLUT_MPORT_76_mask = 1'h1;
  assign cosLUT_MPORT_76_en = reset;
  assign cosLUT_MPORT_77_data = 32'h3f7e3725;
  assign cosLUT_MPORT_77_addr = 11'h4d;
  assign cosLUT_MPORT_77_mask = 1'h1;
  assign cosLUT_MPORT_77_en = reset;
  assign cosLUT_MPORT_78_data = 32'h3f7e2b37;
  assign cosLUT_MPORT_78_addr = 11'h4e;
  assign cosLUT_MPORT_78_mask = 1'h1;
  assign cosLUT_MPORT_78_en = reset;
  assign cosLUT_MPORT_79_data = 32'h3f7e1f22;
  assign cosLUT_MPORT_79_addr = 11'h4f;
  assign cosLUT_MPORT_79_mask = 1'h1;
  assign cosLUT_MPORT_79_en = reset;
  assign cosLUT_MPORT_80_data = 32'h3f7e12e6;
  assign cosLUT_MPORT_80_addr = 11'h50;
  assign cosLUT_MPORT_80_mask = 1'h1;
  assign cosLUT_MPORT_80_en = reset;
  assign cosLUT_MPORT_81_data = 32'h3f7e0682;
  assign cosLUT_MPORT_81_addr = 11'h51;
  assign cosLUT_MPORT_81_mask = 1'h1;
  assign cosLUT_MPORT_81_en = reset;
  assign cosLUT_MPORT_82_data = 32'h3f7df9f8;
  assign cosLUT_MPORT_82_addr = 11'h52;
  assign cosLUT_MPORT_82_mask = 1'h1;
  assign cosLUT_MPORT_82_en = reset;
  assign cosLUT_MPORT_83_data = 32'h3f7ded46;
  assign cosLUT_MPORT_83_addr = 11'h53;
  assign cosLUT_MPORT_83_mask = 1'h1;
  assign cosLUT_MPORT_83_en = reset;
  assign cosLUT_MPORT_84_data = 32'h3f7de06d;
  assign cosLUT_MPORT_84_addr = 11'h54;
  assign cosLUT_MPORT_84_mask = 1'h1;
  assign cosLUT_MPORT_84_en = reset;
  assign cosLUT_MPORT_85_data = 32'h3f7dd36d;
  assign cosLUT_MPORT_85_addr = 11'h55;
  assign cosLUT_MPORT_85_mask = 1'h1;
  assign cosLUT_MPORT_85_en = reset;
  assign cosLUT_MPORT_86_data = 32'h3f7dc645;
  assign cosLUT_MPORT_86_addr = 11'h56;
  assign cosLUT_MPORT_86_mask = 1'h1;
  assign cosLUT_MPORT_86_en = reset;
  assign cosLUT_MPORT_87_data = 32'h3f7db8f7;
  assign cosLUT_MPORT_87_addr = 11'h57;
  assign cosLUT_MPORT_87_mask = 1'h1;
  assign cosLUT_MPORT_87_en = reset;
  assign cosLUT_MPORT_88_data = 32'h3f7dab81;
  assign cosLUT_MPORT_88_addr = 11'h58;
  assign cosLUT_MPORT_88_mask = 1'h1;
  assign cosLUT_MPORT_88_en = reset;
  assign cosLUT_MPORT_89_data = 32'h3f7d9de4;
  assign cosLUT_MPORT_89_addr = 11'h59;
  assign cosLUT_MPORT_89_mask = 1'h1;
  assign cosLUT_MPORT_89_en = reset;
  assign cosLUT_MPORT_90_data = 32'h3f7d9020;
  assign cosLUT_MPORT_90_addr = 11'h5a;
  assign cosLUT_MPORT_90_mask = 1'h1;
  assign cosLUT_MPORT_90_en = reset;
  assign cosLUT_MPORT_91_data = 32'h3f7d8235;
  assign cosLUT_MPORT_91_addr = 11'h5b;
  assign cosLUT_MPORT_91_mask = 1'h1;
  assign cosLUT_MPORT_91_en = reset;
  assign cosLUT_MPORT_92_data = 32'h3f7d7423;
  assign cosLUT_MPORT_92_addr = 11'h5c;
  assign cosLUT_MPORT_92_mask = 1'h1;
  assign cosLUT_MPORT_92_en = reset;
  assign cosLUT_MPORT_93_data = 32'h3f7d65ea;
  assign cosLUT_MPORT_93_addr = 11'h5d;
  assign cosLUT_MPORT_93_mask = 1'h1;
  assign cosLUT_MPORT_93_en = reset;
  assign cosLUT_MPORT_94_data = 32'h3f7d5789;
  assign cosLUT_MPORT_94_addr = 11'h5e;
  assign cosLUT_MPORT_94_mask = 1'h1;
  assign cosLUT_MPORT_94_en = reset;
  assign cosLUT_MPORT_95_data = 32'h3f7d4902;
  assign cosLUT_MPORT_95_addr = 11'h5f;
  assign cosLUT_MPORT_95_mask = 1'h1;
  assign cosLUT_MPORT_95_en = reset;
  assign cosLUT_MPORT_96_data = 32'h3f7d3a53;
  assign cosLUT_MPORT_96_addr = 11'h60;
  assign cosLUT_MPORT_96_mask = 1'h1;
  assign cosLUT_MPORT_96_en = reset;
  assign cosLUT_MPORT_97_data = 32'h3f7d2b7e;
  assign cosLUT_MPORT_97_addr = 11'h61;
  assign cosLUT_MPORT_97_mask = 1'h1;
  assign cosLUT_MPORT_97_en = reset;
  assign cosLUT_MPORT_98_data = 32'h3f7d1c81;
  assign cosLUT_MPORT_98_addr = 11'h62;
  assign cosLUT_MPORT_98_mask = 1'h1;
  assign cosLUT_MPORT_98_en = reset;
  assign cosLUT_MPORT_99_data = 32'h3f7d0d5d;
  assign cosLUT_MPORT_99_addr = 11'h63;
  assign cosLUT_MPORT_99_mask = 1'h1;
  assign cosLUT_MPORT_99_en = reset;
  assign cosLUT_MPORT_100_data = 32'h3f7cfe13;
  assign cosLUT_MPORT_100_addr = 11'h64;
  assign cosLUT_MPORT_100_mask = 1'h1;
  assign cosLUT_MPORT_100_en = reset;
  assign cosLUT_MPORT_101_data = 32'h3f7ceea1;
  assign cosLUT_MPORT_101_addr = 11'h65;
  assign cosLUT_MPORT_101_mask = 1'h1;
  assign cosLUT_MPORT_101_en = reset;
  assign cosLUT_MPORT_102_data = 32'h3f7cdf08;
  assign cosLUT_MPORT_102_addr = 11'h66;
  assign cosLUT_MPORT_102_mask = 1'h1;
  assign cosLUT_MPORT_102_en = reset;
  assign cosLUT_MPORT_103_data = 32'h3f7ccf48;
  assign cosLUT_MPORT_103_addr = 11'h67;
  assign cosLUT_MPORT_103_mask = 1'h1;
  assign cosLUT_MPORT_103_en = reset;
  assign cosLUT_MPORT_104_data = 32'h3f7cbf61;
  assign cosLUT_MPORT_104_addr = 11'h68;
  assign cosLUT_MPORT_104_mask = 1'h1;
  assign cosLUT_MPORT_104_en = reset;
  assign cosLUT_MPORT_105_data = 32'h3f7caf53;
  assign cosLUT_MPORT_105_addr = 11'h69;
  assign cosLUT_MPORT_105_mask = 1'h1;
  assign cosLUT_MPORT_105_en = reset;
  assign cosLUT_MPORT_106_data = 32'h3f7c9f1f;
  assign cosLUT_MPORT_106_addr = 11'h6a;
  assign cosLUT_MPORT_106_mask = 1'h1;
  assign cosLUT_MPORT_106_en = reset;
  assign cosLUT_MPORT_107_data = 32'h3f7c8ec3;
  assign cosLUT_MPORT_107_addr = 11'h6b;
  assign cosLUT_MPORT_107_mask = 1'h1;
  assign cosLUT_MPORT_107_en = reset;
  assign cosLUT_MPORT_108_data = 32'h3f7c7e40;
  assign cosLUT_MPORT_108_addr = 11'h6c;
  assign cosLUT_MPORT_108_mask = 1'h1;
  assign cosLUT_MPORT_108_en = reset;
  assign cosLUT_MPORT_109_data = 32'h3f7c6d96;
  assign cosLUT_MPORT_109_addr = 11'h6d;
  assign cosLUT_MPORT_109_mask = 1'h1;
  assign cosLUT_MPORT_109_en = reset;
  assign cosLUT_MPORT_110_data = 32'h3f7c5cc6;
  assign cosLUT_MPORT_110_addr = 11'h6e;
  assign cosLUT_MPORT_110_mask = 1'h1;
  assign cosLUT_MPORT_110_en = reset;
  assign cosLUT_MPORT_111_data = 32'h3f7c4bce;
  assign cosLUT_MPORT_111_addr = 11'h6f;
  assign cosLUT_MPORT_111_mask = 1'h1;
  assign cosLUT_MPORT_111_en = reset;
  assign cosLUT_MPORT_112_data = 32'h3f7c3aaf;
  assign cosLUT_MPORT_112_addr = 11'h70;
  assign cosLUT_MPORT_112_mask = 1'h1;
  assign cosLUT_MPORT_112_en = reset;
  assign cosLUT_MPORT_113_data = 32'h3f7c296a;
  assign cosLUT_MPORT_113_addr = 11'h71;
  assign cosLUT_MPORT_113_mask = 1'h1;
  assign cosLUT_MPORT_113_en = reset;
  assign cosLUT_MPORT_114_data = 32'h3f7c17fe;
  assign cosLUT_MPORT_114_addr = 11'h72;
  assign cosLUT_MPORT_114_mask = 1'h1;
  assign cosLUT_MPORT_114_en = reset;
  assign cosLUT_MPORT_115_data = 32'h3f7c066a;
  assign cosLUT_MPORT_115_addr = 11'h73;
  assign cosLUT_MPORT_115_mask = 1'h1;
  assign cosLUT_MPORT_115_en = reset;
  assign cosLUT_MPORT_116_data = 32'h3f7bf4b0;
  assign cosLUT_MPORT_116_addr = 11'h74;
  assign cosLUT_MPORT_116_mask = 1'h1;
  assign cosLUT_MPORT_116_en = reset;
  assign cosLUT_MPORT_117_data = 32'h3f7be2cf;
  assign cosLUT_MPORT_117_addr = 11'h75;
  assign cosLUT_MPORT_117_mask = 1'h1;
  assign cosLUT_MPORT_117_en = reset;
  assign cosLUT_MPORT_118_data = 32'h3f7bd0c7;
  assign cosLUT_MPORT_118_addr = 11'h76;
  assign cosLUT_MPORT_118_mask = 1'h1;
  assign cosLUT_MPORT_118_en = reset;
  assign cosLUT_MPORT_119_data = 32'h3f7bbe99;
  assign cosLUT_MPORT_119_addr = 11'h77;
  assign cosLUT_MPORT_119_mask = 1'h1;
  assign cosLUT_MPORT_119_en = reset;
  assign cosLUT_MPORT_120_data = 32'h3f7bac43;
  assign cosLUT_MPORT_120_addr = 11'h78;
  assign cosLUT_MPORT_120_mask = 1'h1;
  assign cosLUT_MPORT_120_en = reset;
  assign cosLUT_MPORT_121_data = 32'h3f7b99c7;
  assign cosLUT_MPORT_121_addr = 11'h79;
  assign cosLUT_MPORT_121_mask = 1'h1;
  assign cosLUT_MPORT_121_en = reset;
  assign cosLUT_MPORT_122_data = 32'h3f7b8723;
  assign cosLUT_MPORT_122_addr = 11'h7a;
  assign cosLUT_MPORT_122_mask = 1'h1;
  assign cosLUT_MPORT_122_en = reset;
  assign cosLUT_MPORT_123_data = 32'h3f7b7459;
  assign cosLUT_MPORT_123_addr = 11'h7b;
  assign cosLUT_MPORT_123_mask = 1'h1;
  assign cosLUT_MPORT_123_en = reset;
  assign cosLUT_MPORT_124_data = 32'h3f7b6169;
  assign cosLUT_MPORT_124_addr = 11'h7c;
  assign cosLUT_MPORT_124_mask = 1'h1;
  assign cosLUT_MPORT_124_en = reset;
  assign cosLUT_MPORT_125_data = 32'h3f7b4e51;
  assign cosLUT_MPORT_125_addr = 11'h7d;
  assign cosLUT_MPORT_125_mask = 1'h1;
  assign cosLUT_MPORT_125_en = reset;
  assign cosLUT_MPORT_126_data = 32'h3f7b3b13;
  assign cosLUT_MPORT_126_addr = 11'h7e;
  assign cosLUT_MPORT_126_mask = 1'h1;
  assign cosLUT_MPORT_126_en = reset;
  assign cosLUT_MPORT_127_data = 32'h3f7b27ad;
  assign cosLUT_MPORT_127_addr = 11'h7f;
  assign cosLUT_MPORT_127_mask = 1'h1;
  assign cosLUT_MPORT_127_en = reset;
  assign cosLUT_MPORT_128_data = 32'h3f7b1422;
  assign cosLUT_MPORT_128_addr = 11'h80;
  assign cosLUT_MPORT_128_mask = 1'h1;
  assign cosLUT_MPORT_128_en = reset;
  assign cosLUT_MPORT_129_data = 32'h3f7b006f;
  assign cosLUT_MPORT_129_addr = 11'h81;
  assign cosLUT_MPORT_129_mask = 1'h1;
  assign cosLUT_MPORT_129_en = reset;
  assign cosLUT_MPORT_130_data = 32'h3f7aec96;
  assign cosLUT_MPORT_130_addr = 11'h82;
  assign cosLUT_MPORT_130_mask = 1'h1;
  assign cosLUT_MPORT_130_en = reset;
  assign cosLUT_MPORT_131_data = 32'h3f7ad895;
  assign cosLUT_MPORT_131_addr = 11'h83;
  assign cosLUT_MPORT_131_mask = 1'h1;
  assign cosLUT_MPORT_131_en = reset;
  assign cosLUT_MPORT_132_data = 32'h3f7ac46f;
  assign cosLUT_MPORT_132_addr = 11'h84;
  assign cosLUT_MPORT_132_mask = 1'h1;
  assign cosLUT_MPORT_132_en = reset;
  assign cosLUT_MPORT_133_data = 32'h3f7ab021;
  assign cosLUT_MPORT_133_addr = 11'h85;
  assign cosLUT_MPORT_133_mask = 1'h1;
  assign cosLUT_MPORT_133_en = reset;
  assign cosLUT_MPORT_134_data = 32'h3f7a9bad;
  assign cosLUT_MPORT_134_addr = 11'h86;
  assign cosLUT_MPORT_134_mask = 1'h1;
  assign cosLUT_MPORT_134_en = reset;
  assign cosLUT_MPORT_135_data = 32'h3f7a8712;
  assign cosLUT_MPORT_135_addr = 11'h87;
  assign cosLUT_MPORT_135_mask = 1'h1;
  assign cosLUT_MPORT_135_en = reset;
  assign cosLUT_MPORT_136_data = 32'h3f7a7251;
  assign cosLUT_MPORT_136_addr = 11'h88;
  assign cosLUT_MPORT_136_mask = 1'h1;
  assign cosLUT_MPORT_136_en = reset;
  assign cosLUT_MPORT_137_data = 32'h3f7a5d69;
  assign cosLUT_MPORT_137_addr = 11'h89;
  assign cosLUT_MPORT_137_mask = 1'h1;
  assign cosLUT_MPORT_137_en = reset;
  assign cosLUT_MPORT_138_data = 32'h3f7a485a;
  assign cosLUT_MPORT_138_addr = 11'h8a;
  assign cosLUT_MPORT_138_mask = 1'h1;
  assign cosLUT_MPORT_138_en = reset;
  assign cosLUT_MPORT_139_data = 32'h3f7a3325;
  assign cosLUT_MPORT_139_addr = 11'h8b;
  assign cosLUT_MPORT_139_mask = 1'h1;
  assign cosLUT_MPORT_139_en = reset;
  assign cosLUT_MPORT_140_data = 32'h3f7a1dc9;
  assign cosLUT_MPORT_140_addr = 11'h8c;
  assign cosLUT_MPORT_140_mask = 1'h1;
  assign cosLUT_MPORT_140_en = reset;
  assign cosLUT_MPORT_141_data = 32'h3f7a0846;
  assign cosLUT_MPORT_141_addr = 11'h8d;
  assign cosLUT_MPORT_141_mask = 1'h1;
  assign cosLUT_MPORT_141_en = reset;
  assign cosLUT_MPORT_142_data = 32'h3f79f29d;
  assign cosLUT_MPORT_142_addr = 11'h8e;
  assign cosLUT_MPORT_142_mask = 1'h1;
  assign cosLUT_MPORT_142_en = reset;
  assign cosLUT_MPORT_143_data = 32'h3f79dccd;
  assign cosLUT_MPORT_143_addr = 11'h8f;
  assign cosLUT_MPORT_143_mask = 1'h1;
  assign cosLUT_MPORT_143_en = reset;
  assign cosLUT_MPORT_144_data = 32'h3f79c6d7;
  assign cosLUT_MPORT_144_addr = 11'h90;
  assign cosLUT_MPORT_144_mask = 1'h1;
  assign cosLUT_MPORT_144_en = reset;
  assign cosLUT_MPORT_145_data = 32'h3f79b0ba;
  assign cosLUT_MPORT_145_addr = 11'h91;
  assign cosLUT_MPORT_145_mask = 1'h1;
  assign cosLUT_MPORT_145_en = reset;
  assign cosLUT_MPORT_146_data = 32'h3f799a77;
  assign cosLUT_MPORT_146_addr = 11'h92;
  assign cosLUT_MPORT_146_mask = 1'h1;
  assign cosLUT_MPORT_146_en = reset;
  assign cosLUT_MPORT_147_data = 32'h3f79840d;
  assign cosLUT_MPORT_147_addr = 11'h93;
  assign cosLUT_MPORT_147_mask = 1'h1;
  assign cosLUT_MPORT_147_en = reset;
  assign cosLUT_MPORT_148_data = 32'h3f796d7d;
  assign cosLUT_MPORT_148_addr = 11'h94;
  assign cosLUT_MPORT_148_mask = 1'h1;
  assign cosLUT_MPORT_148_en = reset;
  assign cosLUT_MPORT_149_data = 32'h3f7956c6;
  assign cosLUT_MPORT_149_addr = 11'h95;
  assign cosLUT_MPORT_149_mask = 1'h1;
  assign cosLUT_MPORT_149_en = reset;
  assign cosLUT_MPORT_150_data = 32'h3f793fe9;
  assign cosLUT_MPORT_150_addr = 11'h96;
  assign cosLUT_MPORT_150_mask = 1'h1;
  assign cosLUT_MPORT_150_en = reset;
  assign cosLUT_MPORT_151_data = 32'h3f7928e5;
  assign cosLUT_MPORT_151_addr = 11'h97;
  assign cosLUT_MPORT_151_mask = 1'h1;
  assign cosLUT_MPORT_151_en = reset;
  assign cosLUT_MPORT_152_data = 32'h3f7911bb;
  assign cosLUT_MPORT_152_addr = 11'h98;
  assign cosLUT_MPORT_152_mask = 1'h1;
  assign cosLUT_MPORT_152_en = reset;
  assign cosLUT_MPORT_153_data = 32'h3f78fa6a;
  assign cosLUT_MPORT_153_addr = 11'h99;
  assign cosLUT_MPORT_153_mask = 1'h1;
  assign cosLUT_MPORT_153_en = reset;
  assign cosLUT_MPORT_154_data = 32'h3f78e2f3;
  assign cosLUT_MPORT_154_addr = 11'h9a;
  assign cosLUT_MPORT_154_mask = 1'h1;
  assign cosLUT_MPORT_154_en = reset;
  assign cosLUT_MPORT_155_data = 32'h3f78cb56;
  assign cosLUT_MPORT_155_addr = 11'h9b;
  assign cosLUT_MPORT_155_mask = 1'h1;
  assign cosLUT_MPORT_155_en = reset;
  assign cosLUT_MPORT_156_data = 32'h3f78b392;
  assign cosLUT_MPORT_156_addr = 11'h9c;
  assign cosLUT_MPORT_156_mask = 1'h1;
  assign cosLUT_MPORT_156_en = reset;
  assign cosLUT_MPORT_157_data = 32'h3f789ba8;
  assign cosLUT_MPORT_157_addr = 11'h9d;
  assign cosLUT_MPORT_157_mask = 1'h1;
  assign cosLUT_MPORT_157_en = reset;
  assign cosLUT_MPORT_158_data = 32'h3f788398;
  assign cosLUT_MPORT_158_addr = 11'h9e;
  assign cosLUT_MPORT_158_mask = 1'h1;
  assign cosLUT_MPORT_158_en = reset;
  assign cosLUT_MPORT_159_data = 32'h3f786b61;
  assign cosLUT_MPORT_159_addr = 11'h9f;
  assign cosLUT_MPORT_159_mask = 1'h1;
  assign cosLUT_MPORT_159_en = reset;
  assign cosLUT_MPORT_160_data = 32'h3f785304;
  assign cosLUT_MPORT_160_addr = 11'ha0;
  assign cosLUT_MPORT_160_mask = 1'h1;
  assign cosLUT_MPORT_160_en = reset;
  assign cosLUT_MPORT_161_data = 32'h3f783a80;
  assign cosLUT_MPORT_161_addr = 11'ha1;
  assign cosLUT_MPORT_161_mask = 1'h1;
  assign cosLUT_MPORT_161_en = reset;
  assign cosLUT_MPORT_162_data = 32'h3f7821d6;
  assign cosLUT_MPORT_162_addr = 11'ha2;
  assign cosLUT_MPORT_162_mask = 1'h1;
  assign cosLUT_MPORT_162_en = reset;
  assign cosLUT_MPORT_163_data = 32'h3f780906;
  assign cosLUT_MPORT_163_addr = 11'ha3;
  assign cosLUT_MPORT_163_mask = 1'h1;
  assign cosLUT_MPORT_163_en = reset;
  assign cosLUT_MPORT_164_data = 32'h3f77f010;
  assign cosLUT_MPORT_164_addr = 11'ha4;
  assign cosLUT_MPORT_164_mask = 1'h1;
  assign cosLUT_MPORT_164_en = reset;
  assign cosLUT_MPORT_165_data = 32'h3f77d6f3;
  assign cosLUT_MPORT_165_addr = 11'ha5;
  assign cosLUT_MPORT_165_mask = 1'h1;
  assign cosLUT_MPORT_165_en = reset;
  assign cosLUT_MPORT_166_data = 32'h3f77bdb0;
  assign cosLUT_MPORT_166_addr = 11'ha6;
  assign cosLUT_MPORT_166_mask = 1'h1;
  assign cosLUT_MPORT_166_en = reset;
  assign cosLUT_MPORT_167_data = 32'h3f77a447;
  assign cosLUT_MPORT_167_addr = 11'ha7;
  assign cosLUT_MPORT_167_mask = 1'h1;
  assign cosLUT_MPORT_167_en = reset;
  assign cosLUT_MPORT_168_data = 32'h3f778ab8;
  assign cosLUT_MPORT_168_addr = 11'ha8;
  assign cosLUT_MPORT_168_mask = 1'h1;
  assign cosLUT_MPORT_168_en = reset;
  assign cosLUT_MPORT_169_data = 32'h3f777103;
  assign cosLUT_MPORT_169_addr = 11'ha9;
  assign cosLUT_MPORT_169_mask = 1'h1;
  assign cosLUT_MPORT_169_en = reset;
  assign cosLUT_MPORT_170_data = 32'h3f775727;
  assign cosLUT_MPORT_170_addr = 11'haa;
  assign cosLUT_MPORT_170_mask = 1'h1;
  assign cosLUT_MPORT_170_en = reset;
  assign cosLUT_MPORT_171_data = 32'h3f773d25;
  assign cosLUT_MPORT_171_addr = 11'hab;
  assign cosLUT_MPORT_171_mask = 1'h1;
  assign cosLUT_MPORT_171_en = reset;
  assign cosLUT_MPORT_172_data = 32'h3f7722fd;
  assign cosLUT_MPORT_172_addr = 11'hac;
  assign cosLUT_MPORT_172_mask = 1'h1;
  assign cosLUT_MPORT_172_en = reset;
  assign cosLUT_MPORT_173_data = 32'h3f7708af;
  assign cosLUT_MPORT_173_addr = 11'had;
  assign cosLUT_MPORT_173_mask = 1'h1;
  assign cosLUT_MPORT_173_en = reset;
  assign cosLUT_MPORT_174_data = 32'h3f76ee3b;
  assign cosLUT_MPORT_174_addr = 11'hae;
  assign cosLUT_MPORT_174_mask = 1'h1;
  assign cosLUT_MPORT_174_en = reset;
  assign cosLUT_MPORT_175_data = 32'h3f76d3a1;
  assign cosLUT_MPORT_175_addr = 11'haf;
  assign cosLUT_MPORT_175_mask = 1'h1;
  assign cosLUT_MPORT_175_en = reset;
  assign cosLUT_MPORT_176_data = 32'h3f76b8e0;
  assign cosLUT_MPORT_176_addr = 11'hb0;
  assign cosLUT_MPORT_176_mask = 1'h1;
  assign cosLUT_MPORT_176_en = reset;
  assign cosLUT_MPORT_177_data = 32'h3f769dfa;
  assign cosLUT_MPORT_177_addr = 11'hb1;
  assign cosLUT_MPORT_177_mask = 1'h1;
  assign cosLUT_MPORT_177_en = reset;
  assign cosLUT_MPORT_178_data = 32'h3f7682ed;
  assign cosLUT_MPORT_178_addr = 11'hb2;
  assign cosLUT_MPORT_178_mask = 1'h1;
  assign cosLUT_MPORT_178_en = reset;
  assign cosLUT_MPORT_179_data = 32'h3f7667bb;
  assign cosLUT_MPORT_179_addr = 11'hb3;
  assign cosLUT_MPORT_179_mask = 1'h1;
  assign cosLUT_MPORT_179_en = reset;
  assign cosLUT_MPORT_180_data = 32'h3f764c62;
  assign cosLUT_MPORT_180_addr = 11'hb4;
  assign cosLUT_MPORT_180_mask = 1'h1;
  assign cosLUT_MPORT_180_en = reset;
  assign cosLUT_MPORT_181_data = 32'h3f7630e4;
  assign cosLUT_MPORT_181_addr = 11'hb5;
  assign cosLUT_MPORT_181_mask = 1'h1;
  assign cosLUT_MPORT_181_en = reset;
  assign cosLUT_MPORT_182_data = 32'h3f76153f;
  assign cosLUT_MPORT_182_addr = 11'hb6;
  assign cosLUT_MPORT_182_mask = 1'h1;
  assign cosLUT_MPORT_182_en = reset;
  assign cosLUT_MPORT_183_data = 32'h3f75f975;
  assign cosLUT_MPORT_183_addr = 11'hb7;
  assign cosLUT_MPORT_183_mask = 1'h1;
  assign cosLUT_MPORT_183_en = reset;
  assign cosLUT_MPORT_184_data = 32'h3f75dd84;
  assign cosLUT_MPORT_184_addr = 11'hb8;
  assign cosLUT_MPORT_184_mask = 1'h1;
  assign cosLUT_MPORT_184_en = reset;
  assign cosLUT_MPORT_185_data = 32'h3f75c16e;
  assign cosLUT_MPORT_185_addr = 11'hb9;
  assign cosLUT_MPORT_185_mask = 1'h1;
  assign cosLUT_MPORT_185_en = reset;
  assign cosLUT_MPORT_186_data = 32'h3f75a531;
  assign cosLUT_MPORT_186_addr = 11'hba;
  assign cosLUT_MPORT_186_mask = 1'h1;
  assign cosLUT_MPORT_186_en = reset;
  assign cosLUT_MPORT_187_data = 32'h3f7588cf;
  assign cosLUT_MPORT_187_addr = 11'hbb;
  assign cosLUT_MPORT_187_mask = 1'h1;
  assign cosLUT_MPORT_187_en = reset;
  assign cosLUT_MPORT_188_data = 32'h3f756c47;
  assign cosLUT_MPORT_188_addr = 11'hbc;
  assign cosLUT_MPORT_188_mask = 1'h1;
  assign cosLUT_MPORT_188_en = reset;
  assign cosLUT_MPORT_189_data = 32'h3f754f99;
  assign cosLUT_MPORT_189_addr = 11'hbd;
  assign cosLUT_MPORT_189_mask = 1'h1;
  assign cosLUT_MPORT_189_en = reset;
  assign cosLUT_MPORT_190_data = 32'h3f7532c5;
  assign cosLUT_MPORT_190_addr = 11'hbe;
  assign cosLUT_MPORT_190_mask = 1'h1;
  assign cosLUT_MPORT_190_en = reset;
  assign cosLUT_MPORT_191_data = 32'h3f7515cc;
  assign cosLUT_MPORT_191_addr = 11'hbf;
  assign cosLUT_MPORT_191_mask = 1'h1;
  assign cosLUT_MPORT_191_en = reset;
  assign cosLUT_MPORT_192_data = 32'h3f74f8ac;
  assign cosLUT_MPORT_192_addr = 11'hc0;
  assign cosLUT_MPORT_192_mask = 1'h1;
  assign cosLUT_MPORT_192_en = reset;
  assign cosLUT_MPORT_193_data = 32'h3f74db67;
  assign cosLUT_MPORT_193_addr = 11'hc1;
  assign cosLUT_MPORT_193_mask = 1'h1;
  assign cosLUT_MPORT_193_en = reset;
  assign cosLUT_MPORT_194_data = 32'h3f74bdfc;
  assign cosLUT_MPORT_194_addr = 11'hc2;
  assign cosLUT_MPORT_194_mask = 1'h1;
  assign cosLUT_MPORT_194_en = reset;
  assign cosLUT_MPORT_195_data = 32'h3f74a06b;
  assign cosLUT_MPORT_195_addr = 11'hc3;
  assign cosLUT_MPORT_195_mask = 1'h1;
  assign cosLUT_MPORT_195_en = reset;
  assign cosLUT_MPORT_196_data = 32'h3f7482b5;
  assign cosLUT_MPORT_196_addr = 11'hc4;
  assign cosLUT_MPORT_196_mask = 1'h1;
  assign cosLUT_MPORT_196_en = reset;
  assign cosLUT_MPORT_197_data = 32'h3f7464d9;
  assign cosLUT_MPORT_197_addr = 11'hc5;
  assign cosLUT_MPORT_197_mask = 1'h1;
  assign cosLUT_MPORT_197_en = reset;
  assign cosLUT_MPORT_198_data = 32'h3f7446d7;
  assign cosLUT_MPORT_198_addr = 11'hc6;
  assign cosLUT_MPORT_198_mask = 1'h1;
  assign cosLUT_MPORT_198_en = reset;
  assign cosLUT_MPORT_199_data = 32'h3f7428af;
  assign cosLUT_MPORT_199_addr = 11'hc7;
  assign cosLUT_MPORT_199_mask = 1'h1;
  assign cosLUT_MPORT_199_en = reset;
  assign cosLUT_MPORT_200_data = 32'h3f740a62;
  assign cosLUT_MPORT_200_addr = 11'hc8;
  assign cosLUT_MPORT_200_mask = 1'h1;
  assign cosLUT_MPORT_200_en = reset;
  assign cosLUT_MPORT_201_data = 32'h3f73ebef;
  assign cosLUT_MPORT_201_addr = 11'hc9;
  assign cosLUT_MPORT_201_mask = 1'h1;
  assign cosLUT_MPORT_201_en = reset;
  assign cosLUT_MPORT_202_data = 32'h3f73cd56;
  assign cosLUT_MPORT_202_addr = 11'hca;
  assign cosLUT_MPORT_202_mask = 1'h1;
  assign cosLUT_MPORT_202_en = reset;
  assign cosLUT_MPORT_203_data = 32'h3f73ae98;
  assign cosLUT_MPORT_203_addr = 11'hcb;
  assign cosLUT_MPORT_203_mask = 1'h1;
  assign cosLUT_MPORT_203_en = reset;
  assign cosLUT_MPORT_204_data = 32'h3f738fb4;
  assign cosLUT_MPORT_204_addr = 11'hcc;
  assign cosLUT_MPORT_204_mask = 1'h1;
  assign cosLUT_MPORT_204_en = reset;
  assign cosLUT_MPORT_205_data = 32'h3f7370ab;
  assign cosLUT_MPORT_205_addr = 11'hcd;
  assign cosLUT_MPORT_205_mask = 1'h1;
  assign cosLUT_MPORT_205_en = reset;
  assign cosLUT_MPORT_206_data = 32'h3f73517c;
  assign cosLUT_MPORT_206_addr = 11'hce;
  assign cosLUT_MPORT_206_mask = 1'h1;
  assign cosLUT_MPORT_206_en = reset;
  assign cosLUT_MPORT_207_data = 32'h3f733227;
  assign cosLUT_MPORT_207_addr = 11'hcf;
  assign cosLUT_MPORT_207_mask = 1'h1;
  assign cosLUT_MPORT_207_en = reset;
  assign cosLUT_MPORT_208_data = 32'h3f7312ad;
  assign cosLUT_MPORT_208_addr = 11'hd0;
  assign cosLUT_MPORT_208_mask = 1'h1;
  assign cosLUT_MPORT_208_en = reset;
  assign cosLUT_MPORT_209_data = 32'h3f72f30e;
  assign cosLUT_MPORT_209_addr = 11'hd1;
  assign cosLUT_MPORT_209_mask = 1'h1;
  assign cosLUT_MPORT_209_en = reset;
  assign cosLUT_MPORT_210_data = 32'h3f72d349;
  assign cosLUT_MPORT_210_addr = 11'hd2;
  assign cosLUT_MPORT_210_mask = 1'h1;
  assign cosLUT_MPORT_210_en = reset;
  assign cosLUT_MPORT_211_data = 32'h3f72b35e;
  assign cosLUT_MPORT_211_addr = 11'hd3;
  assign cosLUT_MPORT_211_mask = 1'h1;
  assign cosLUT_MPORT_211_en = reset;
  assign cosLUT_MPORT_212_data = 32'h3f72934e;
  assign cosLUT_MPORT_212_addr = 11'hd4;
  assign cosLUT_MPORT_212_mask = 1'h1;
  assign cosLUT_MPORT_212_en = reset;
  assign cosLUT_MPORT_213_data = 32'h3f727319;
  assign cosLUT_MPORT_213_addr = 11'hd5;
  assign cosLUT_MPORT_213_mask = 1'h1;
  assign cosLUT_MPORT_213_en = reset;
  assign cosLUT_MPORT_214_data = 32'h3f7252be;
  assign cosLUT_MPORT_214_addr = 11'hd6;
  assign cosLUT_MPORT_214_mask = 1'h1;
  assign cosLUT_MPORT_214_en = reset;
  assign cosLUT_MPORT_215_data = 32'h3f72323e;
  assign cosLUT_MPORT_215_addr = 11'hd7;
  assign cosLUT_MPORT_215_mask = 1'h1;
  assign cosLUT_MPORT_215_en = reset;
  assign cosLUT_MPORT_216_data = 32'h3f721199;
  assign cosLUT_MPORT_216_addr = 11'hd8;
  assign cosLUT_MPORT_216_mask = 1'h1;
  assign cosLUT_MPORT_216_en = reset;
  assign cosLUT_MPORT_217_data = 32'h3f71f0ce;
  assign cosLUT_MPORT_217_addr = 11'hd9;
  assign cosLUT_MPORT_217_mask = 1'h1;
  assign cosLUT_MPORT_217_en = reset;
  assign cosLUT_MPORT_218_data = 32'h3f71cfde;
  assign cosLUT_MPORT_218_addr = 11'hda;
  assign cosLUT_MPORT_218_mask = 1'h1;
  assign cosLUT_MPORT_218_en = reset;
  assign cosLUT_MPORT_219_data = 32'h3f71aec8;
  assign cosLUT_MPORT_219_addr = 11'hdb;
  assign cosLUT_MPORT_219_mask = 1'h1;
  assign cosLUT_MPORT_219_en = reset;
  assign cosLUT_MPORT_220_data = 32'h3f718d8d;
  assign cosLUT_MPORT_220_addr = 11'hdc;
  assign cosLUT_MPORT_220_mask = 1'h1;
  assign cosLUT_MPORT_220_en = reset;
  assign cosLUT_MPORT_221_data = 32'h3f716c2d;
  assign cosLUT_MPORT_221_addr = 11'hdd;
  assign cosLUT_MPORT_221_mask = 1'h1;
  assign cosLUT_MPORT_221_en = reset;
  assign cosLUT_MPORT_222_data = 32'h3f714aa8;
  assign cosLUT_MPORT_222_addr = 11'hde;
  assign cosLUT_MPORT_222_mask = 1'h1;
  assign cosLUT_MPORT_222_en = reset;
  assign cosLUT_MPORT_223_data = 32'h3f7128fe;
  assign cosLUT_MPORT_223_addr = 11'hdf;
  assign cosLUT_MPORT_223_mask = 1'h1;
  assign cosLUT_MPORT_223_en = reset;
  assign cosLUT_MPORT_224_data = 32'h3f71072e;
  assign cosLUT_MPORT_224_addr = 11'he0;
  assign cosLUT_MPORT_224_mask = 1'h1;
  assign cosLUT_MPORT_224_en = reset;
  assign cosLUT_MPORT_225_data = 32'h3f70e539;
  assign cosLUT_MPORT_225_addr = 11'he1;
  assign cosLUT_MPORT_225_mask = 1'h1;
  assign cosLUT_MPORT_225_en = reset;
  assign cosLUT_MPORT_226_data = 32'h3f70c31f;
  assign cosLUT_MPORT_226_addr = 11'he2;
  assign cosLUT_MPORT_226_mask = 1'h1;
  assign cosLUT_MPORT_226_en = reset;
  assign cosLUT_MPORT_227_data = 32'h3f70a0e0;
  assign cosLUT_MPORT_227_addr = 11'he3;
  assign cosLUT_MPORT_227_mask = 1'h1;
  assign cosLUT_MPORT_227_en = reset;
  assign cosLUT_MPORT_228_data = 32'h3f707e7b;
  assign cosLUT_MPORT_228_addr = 11'he4;
  assign cosLUT_MPORT_228_mask = 1'h1;
  assign cosLUT_MPORT_228_en = reset;
  assign cosLUT_MPORT_229_data = 32'h3f705bf2;
  assign cosLUT_MPORT_229_addr = 11'he5;
  assign cosLUT_MPORT_229_mask = 1'h1;
  assign cosLUT_MPORT_229_en = reset;
  assign cosLUT_MPORT_230_data = 32'h3f703943;
  assign cosLUT_MPORT_230_addr = 11'he6;
  assign cosLUT_MPORT_230_mask = 1'h1;
  assign cosLUT_MPORT_230_en = reset;
  assign cosLUT_MPORT_231_data = 32'h3f701670;
  assign cosLUT_MPORT_231_addr = 11'he7;
  assign cosLUT_MPORT_231_mask = 1'h1;
  assign cosLUT_MPORT_231_en = reset;
  assign cosLUT_MPORT_232_data = 32'h3f6ff377;
  assign cosLUT_MPORT_232_addr = 11'he8;
  assign cosLUT_MPORT_232_mask = 1'h1;
  assign cosLUT_MPORT_232_en = reset;
  assign cosLUT_MPORT_233_data = 32'h3f6fd059;
  assign cosLUT_MPORT_233_addr = 11'he9;
  assign cosLUT_MPORT_233_mask = 1'h1;
  assign cosLUT_MPORT_233_en = reset;
  assign cosLUT_MPORT_234_data = 32'h3f6fad17;
  assign cosLUT_MPORT_234_addr = 11'hea;
  assign cosLUT_MPORT_234_mask = 1'h1;
  assign cosLUT_MPORT_234_en = reset;
  assign cosLUT_MPORT_235_data = 32'h3f6f89af;
  assign cosLUT_MPORT_235_addr = 11'heb;
  assign cosLUT_MPORT_235_mask = 1'h1;
  assign cosLUT_MPORT_235_en = reset;
  assign cosLUT_MPORT_236_data = 32'h3f6f6622;
  assign cosLUT_MPORT_236_addr = 11'hec;
  assign cosLUT_MPORT_236_mask = 1'h1;
  assign cosLUT_MPORT_236_en = reset;
  assign cosLUT_MPORT_237_data = 32'h3f6f4271;
  assign cosLUT_MPORT_237_addr = 11'hed;
  assign cosLUT_MPORT_237_mask = 1'h1;
  assign cosLUT_MPORT_237_en = reset;
  assign cosLUT_MPORT_238_data = 32'h3f6f1e9a;
  assign cosLUT_MPORT_238_addr = 11'hee;
  assign cosLUT_MPORT_238_mask = 1'h1;
  assign cosLUT_MPORT_238_en = reset;
  assign cosLUT_MPORT_239_data = 32'h3f6efa9f;
  assign cosLUT_MPORT_239_addr = 11'hef;
  assign cosLUT_MPORT_239_mask = 1'h1;
  assign cosLUT_MPORT_239_en = reset;
  assign cosLUT_MPORT_240_data = 32'h3f6ed67f;
  assign cosLUT_MPORT_240_addr = 11'hf0;
  assign cosLUT_MPORT_240_mask = 1'h1;
  assign cosLUT_MPORT_240_en = reset;
  assign cosLUT_MPORT_241_data = 32'h3f6eb23a;
  assign cosLUT_MPORT_241_addr = 11'hf1;
  assign cosLUT_MPORT_241_mask = 1'h1;
  assign cosLUT_MPORT_241_en = reset;
  assign cosLUT_MPORT_242_data = 32'h3f6e8dd0;
  assign cosLUT_MPORT_242_addr = 11'hf2;
  assign cosLUT_MPORT_242_mask = 1'h1;
  assign cosLUT_MPORT_242_en = reset;
  assign cosLUT_MPORT_243_data = 32'h3f6e6941;
  assign cosLUT_MPORT_243_addr = 11'hf3;
  assign cosLUT_MPORT_243_mask = 1'h1;
  assign cosLUT_MPORT_243_en = reset;
  assign cosLUT_MPORT_244_data = 32'h3f6e448e;
  assign cosLUT_MPORT_244_addr = 11'hf4;
  assign cosLUT_MPORT_244_mask = 1'h1;
  assign cosLUT_MPORT_244_en = reset;
  assign cosLUT_MPORT_245_data = 32'h3f6e1fb5;
  assign cosLUT_MPORT_245_addr = 11'hf5;
  assign cosLUT_MPORT_245_mask = 1'h1;
  assign cosLUT_MPORT_245_en = reset;
  assign cosLUT_MPORT_246_data = 32'h3f6dfab8;
  assign cosLUT_MPORT_246_addr = 11'hf6;
  assign cosLUT_MPORT_246_mask = 1'h1;
  assign cosLUT_MPORT_246_en = reset;
  assign cosLUT_MPORT_247_data = 32'h3f6dd597;
  assign cosLUT_MPORT_247_addr = 11'hf7;
  assign cosLUT_MPORT_247_mask = 1'h1;
  assign cosLUT_MPORT_247_en = reset;
  assign cosLUT_MPORT_248_data = 32'h3f6db050;
  assign cosLUT_MPORT_248_addr = 11'hf8;
  assign cosLUT_MPORT_248_mask = 1'h1;
  assign cosLUT_MPORT_248_en = reset;
  assign cosLUT_MPORT_249_data = 32'h3f6d8ae5;
  assign cosLUT_MPORT_249_addr = 11'hf9;
  assign cosLUT_MPORT_249_mask = 1'h1;
  assign cosLUT_MPORT_249_en = reset;
  assign cosLUT_MPORT_250_data = 32'h3f6d6555;
  assign cosLUT_MPORT_250_addr = 11'hfa;
  assign cosLUT_MPORT_250_mask = 1'h1;
  assign cosLUT_MPORT_250_en = reset;
  assign cosLUT_MPORT_251_data = 32'h3f6d3fa1;
  assign cosLUT_MPORT_251_addr = 11'hfb;
  assign cosLUT_MPORT_251_mask = 1'h1;
  assign cosLUT_MPORT_251_en = reset;
  assign cosLUT_MPORT_252_data = 32'h3f6d19c8;
  assign cosLUT_MPORT_252_addr = 11'hfc;
  assign cosLUT_MPORT_252_mask = 1'h1;
  assign cosLUT_MPORT_252_en = reset;
  assign cosLUT_MPORT_253_data = 32'h3f6cf3cb;
  assign cosLUT_MPORT_253_addr = 11'hfd;
  assign cosLUT_MPORT_253_mask = 1'h1;
  assign cosLUT_MPORT_253_en = reset;
  assign cosLUT_MPORT_254_data = 32'h3f6ccda8;
  assign cosLUT_MPORT_254_addr = 11'hfe;
  assign cosLUT_MPORT_254_mask = 1'h1;
  assign cosLUT_MPORT_254_en = reset;
  assign cosLUT_MPORT_255_data = 32'h3f6ca762;
  assign cosLUT_MPORT_255_addr = 11'hff;
  assign cosLUT_MPORT_255_mask = 1'h1;
  assign cosLUT_MPORT_255_en = reset;
  assign cosLUT_MPORT_256_data = 32'h3f6c80f7;
  assign cosLUT_MPORT_256_addr = 11'h100;
  assign cosLUT_MPORT_256_mask = 1'h1;
  assign cosLUT_MPORT_256_en = reset;
  assign cosLUT_MPORT_257_data = 32'h3f6c5a67;
  assign cosLUT_MPORT_257_addr = 11'h101;
  assign cosLUT_MPORT_257_mask = 1'h1;
  assign cosLUT_MPORT_257_en = reset;
  assign cosLUT_MPORT_258_data = 32'h3f6c33b3;
  assign cosLUT_MPORT_258_addr = 11'h102;
  assign cosLUT_MPORT_258_mask = 1'h1;
  assign cosLUT_MPORT_258_en = reset;
  assign cosLUT_MPORT_259_data = 32'h3f6c0cda;
  assign cosLUT_MPORT_259_addr = 11'h103;
  assign cosLUT_MPORT_259_mask = 1'h1;
  assign cosLUT_MPORT_259_en = reset;
  assign cosLUT_MPORT_260_data = 32'h3f6be5dd;
  assign cosLUT_MPORT_260_addr = 11'h104;
  assign cosLUT_MPORT_260_mask = 1'h1;
  assign cosLUT_MPORT_260_en = reset;
  assign cosLUT_MPORT_261_data = 32'h3f6bbebc;
  assign cosLUT_MPORT_261_addr = 11'h105;
  assign cosLUT_MPORT_261_mask = 1'h1;
  assign cosLUT_MPORT_261_en = reset;
  assign cosLUT_MPORT_262_data = 32'h3f6b9776;
  assign cosLUT_MPORT_262_addr = 11'h106;
  assign cosLUT_MPORT_262_mask = 1'h1;
  assign cosLUT_MPORT_262_en = reset;
  assign cosLUT_MPORT_263_data = 32'h3f6b700c;
  assign cosLUT_MPORT_263_addr = 11'h107;
  assign cosLUT_MPORT_263_mask = 1'h1;
  assign cosLUT_MPORT_263_en = reset;
  assign cosLUT_MPORT_264_data = 32'h3f6b487e;
  assign cosLUT_MPORT_264_addr = 11'h108;
  assign cosLUT_MPORT_264_mask = 1'h1;
  assign cosLUT_MPORT_264_en = reset;
  assign cosLUT_MPORT_265_data = 32'h3f6b20cb;
  assign cosLUT_MPORT_265_addr = 11'h109;
  assign cosLUT_MPORT_265_mask = 1'h1;
  assign cosLUT_MPORT_265_en = reset;
  assign cosLUT_MPORT_266_data = 32'h3f6af8f4;
  assign cosLUT_MPORT_266_addr = 11'h10a;
  assign cosLUT_MPORT_266_mask = 1'h1;
  assign cosLUT_MPORT_266_en = reset;
  assign cosLUT_MPORT_267_data = 32'h3f6ad0f9;
  assign cosLUT_MPORT_267_addr = 11'h10b;
  assign cosLUT_MPORT_267_mask = 1'h1;
  assign cosLUT_MPORT_267_en = reset;
  assign cosLUT_MPORT_268_data = 32'h3f6aa8d9;
  assign cosLUT_MPORT_268_addr = 11'h10c;
  assign cosLUT_MPORT_268_mask = 1'h1;
  assign cosLUT_MPORT_268_en = reset;
  assign cosLUT_MPORT_269_data = 32'h3f6a8096;
  assign cosLUT_MPORT_269_addr = 11'h10d;
  assign cosLUT_MPORT_269_mask = 1'h1;
  assign cosLUT_MPORT_269_en = reset;
  assign cosLUT_MPORT_270_data = 32'h3f6a582e;
  assign cosLUT_MPORT_270_addr = 11'h10e;
  assign cosLUT_MPORT_270_mask = 1'h1;
  assign cosLUT_MPORT_270_en = reset;
  assign cosLUT_MPORT_271_data = 32'h3f6a2fa2;
  assign cosLUT_MPORT_271_addr = 11'h10f;
  assign cosLUT_MPORT_271_mask = 1'h1;
  assign cosLUT_MPORT_271_en = reset;
  assign cosLUT_MPORT_272_data = 32'h3f6a06f2;
  assign cosLUT_MPORT_272_addr = 11'h110;
  assign cosLUT_MPORT_272_mask = 1'h1;
  assign cosLUT_MPORT_272_en = reset;
  assign cosLUT_MPORT_273_data = 32'h3f69de1d;
  assign cosLUT_MPORT_273_addr = 11'h111;
  assign cosLUT_MPORT_273_mask = 1'h1;
  assign cosLUT_MPORT_273_en = reset;
  assign cosLUT_MPORT_274_data = 32'h3f69b525;
  assign cosLUT_MPORT_274_addr = 11'h112;
  assign cosLUT_MPORT_274_mask = 1'h1;
  assign cosLUT_MPORT_274_en = reset;
  assign cosLUT_MPORT_275_data = 32'h3f698c09;
  assign cosLUT_MPORT_275_addr = 11'h113;
  assign cosLUT_MPORT_275_mask = 1'h1;
  assign cosLUT_MPORT_275_en = reset;
  assign cosLUT_MPORT_276_data = 32'h3f6962c8;
  assign cosLUT_MPORT_276_addr = 11'h114;
  assign cosLUT_MPORT_276_mask = 1'h1;
  assign cosLUT_MPORT_276_en = reset;
  assign cosLUT_MPORT_277_data = 32'h3f693964;
  assign cosLUT_MPORT_277_addr = 11'h115;
  assign cosLUT_MPORT_277_mask = 1'h1;
  assign cosLUT_MPORT_277_en = reset;
  assign cosLUT_MPORT_278_data = 32'h3f690fdb;
  assign cosLUT_MPORT_278_addr = 11'h116;
  assign cosLUT_MPORT_278_mask = 1'h1;
  assign cosLUT_MPORT_278_en = reset;
  assign cosLUT_MPORT_279_data = 32'h3f68e62f;
  assign cosLUT_MPORT_279_addr = 11'h117;
  assign cosLUT_MPORT_279_mask = 1'h1;
  assign cosLUT_MPORT_279_en = reset;
  assign cosLUT_MPORT_280_data = 32'h3f68bc5f;
  assign cosLUT_MPORT_280_addr = 11'h118;
  assign cosLUT_MPORT_280_mask = 1'h1;
  assign cosLUT_MPORT_280_en = reset;
  assign cosLUT_MPORT_281_data = 32'h3f68926b;
  assign cosLUT_MPORT_281_addr = 11'h119;
  assign cosLUT_MPORT_281_mask = 1'h1;
  assign cosLUT_MPORT_281_en = reset;
  assign cosLUT_MPORT_282_data = 32'h3f686852;
  assign cosLUT_MPORT_282_addr = 11'h11a;
  assign cosLUT_MPORT_282_mask = 1'h1;
  assign cosLUT_MPORT_282_en = reset;
  assign cosLUT_MPORT_283_data = 32'h3f683e16;
  assign cosLUT_MPORT_283_addr = 11'h11b;
  assign cosLUT_MPORT_283_mask = 1'h1;
  assign cosLUT_MPORT_283_en = reset;
  assign cosLUT_MPORT_284_data = 32'h3f6813b7;
  assign cosLUT_MPORT_284_addr = 11'h11c;
  assign cosLUT_MPORT_284_mask = 1'h1;
  assign cosLUT_MPORT_284_en = reset;
  assign cosLUT_MPORT_285_data = 32'h3f67e933;
  assign cosLUT_MPORT_285_addr = 11'h11d;
  assign cosLUT_MPORT_285_mask = 1'h1;
  assign cosLUT_MPORT_285_en = reset;
  assign cosLUT_MPORT_286_data = 32'h3f67be8c;
  assign cosLUT_MPORT_286_addr = 11'h11e;
  assign cosLUT_MPORT_286_mask = 1'h1;
  assign cosLUT_MPORT_286_en = reset;
  assign cosLUT_MPORT_287_data = 32'h3f6793c1;
  assign cosLUT_MPORT_287_addr = 11'h11f;
  assign cosLUT_MPORT_287_mask = 1'h1;
  assign cosLUT_MPORT_287_en = reset;
  assign cosLUT_MPORT_288_data = 32'h3f6768d2;
  assign cosLUT_MPORT_288_addr = 11'h120;
  assign cosLUT_MPORT_288_mask = 1'h1;
  assign cosLUT_MPORT_288_en = reset;
  assign cosLUT_MPORT_289_data = 32'h3f673dbf;
  assign cosLUT_MPORT_289_addr = 11'h121;
  assign cosLUT_MPORT_289_mask = 1'h1;
  assign cosLUT_MPORT_289_en = reset;
  assign cosLUT_MPORT_290_data = 32'h3f671289;
  assign cosLUT_MPORT_290_addr = 11'h122;
  assign cosLUT_MPORT_290_mask = 1'h1;
  assign cosLUT_MPORT_290_en = reset;
  assign cosLUT_MPORT_291_data = 32'h3f66e72f;
  assign cosLUT_MPORT_291_addr = 11'h123;
  assign cosLUT_MPORT_291_mask = 1'h1;
  assign cosLUT_MPORT_291_en = reset;
  assign cosLUT_MPORT_292_data = 32'h3f66bbb1;
  assign cosLUT_MPORT_292_addr = 11'h124;
  assign cosLUT_MPORT_292_mask = 1'h1;
  assign cosLUT_MPORT_292_en = reset;
  assign cosLUT_MPORT_293_data = 32'h3f669010;
  assign cosLUT_MPORT_293_addr = 11'h125;
  assign cosLUT_MPORT_293_mask = 1'h1;
  assign cosLUT_MPORT_293_en = reset;
  assign cosLUT_MPORT_294_data = 32'h3f66644c;
  assign cosLUT_MPORT_294_addr = 11'h126;
  assign cosLUT_MPORT_294_mask = 1'h1;
  assign cosLUT_MPORT_294_en = reset;
  assign cosLUT_MPORT_295_data = 32'h3f663863;
  assign cosLUT_MPORT_295_addr = 11'h127;
  assign cosLUT_MPORT_295_mask = 1'h1;
  assign cosLUT_MPORT_295_en = reset;
  assign cosLUT_MPORT_296_data = 32'h3f660c58;
  assign cosLUT_MPORT_296_addr = 11'h128;
  assign cosLUT_MPORT_296_mask = 1'h1;
  assign cosLUT_MPORT_296_en = reset;
  assign cosLUT_MPORT_297_data = 32'h3f65e028;
  assign cosLUT_MPORT_297_addr = 11'h129;
  assign cosLUT_MPORT_297_mask = 1'h1;
  assign cosLUT_MPORT_297_en = reset;
  assign cosLUT_MPORT_298_data = 32'h3f65b3d6;
  assign cosLUT_MPORT_298_addr = 11'h12a;
  assign cosLUT_MPORT_298_mask = 1'h1;
  assign cosLUT_MPORT_298_en = reset;
  assign cosLUT_MPORT_299_data = 32'h3f65875f;
  assign cosLUT_MPORT_299_addr = 11'h12b;
  assign cosLUT_MPORT_299_mask = 1'h1;
  assign cosLUT_MPORT_299_en = reset;
  assign cosLUT_MPORT_300_data = 32'h3f655ac6;
  assign cosLUT_MPORT_300_addr = 11'h12c;
  assign cosLUT_MPORT_300_mask = 1'h1;
  assign cosLUT_MPORT_300_en = reset;
  assign cosLUT_MPORT_301_data = 32'h3f652e09;
  assign cosLUT_MPORT_301_addr = 11'h12d;
  assign cosLUT_MPORT_301_mask = 1'h1;
  assign cosLUT_MPORT_301_en = reset;
  assign cosLUT_MPORT_302_data = 32'h3f650129;
  assign cosLUT_MPORT_302_addr = 11'h12e;
  assign cosLUT_MPORT_302_mask = 1'h1;
  assign cosLUT_MPORT_302_en = reset;
  assign cosLUT_MPORT_303_data = 32'h3f64d425;
  assign cosLUT_MPORT_303_addr = 11'h12f;
  assign cosLUT_MPORT_303_mask = 1'h1;
  assign cosLUT_MPORT_303_en = reset;
  assign cosLUT_MPORT_304_data = 32'h3f64a6fe;
  assign cosLUT_MPORT_304_addr = 11'h130;
  assign cosLUT_MPORT_304_mask = 1'h1;
  assign cosLUT_MPORT_304_en = reset;
  assign cosLUT_MPORT_305_data = 32'h3f6479b4;
  assign cosLUT_MPORT_305_addr = 11'h131;
  assign cosLUT_MPORT_305_mask = 1'h1;
  assign cosLUT_MPORT_305_en = reset;
  assign cosLUT_MPORT_306_data = 32'h3f644c46;
  assign cosLUT_MPORT_306_addr = 11'h132;
  assign cosLUT_MPORT_306_mask = 1'h1;
  assign cosLUT_MPORT_306_en = reset;
  assign cosLUT_MPORT_307_data = 32'h3f641eb5;
  assign cosLUT_MPORT_307_addr = 11'h133;
  assign cosLUT_MPORT_307_mask = 1'h1;
  assign cosLUT_MPORT_307_en = reset;
  assign cosLUT_MPORT_308_data = 32'h3f63f102;
  assign cosLUT_MPORT_308_addr = 11'h134;
  assign cosLUT_MPORT_308_mask = 1'h1;
  assign cosLUT_MPORT_308_en = reset;
  assign cosLUT_MPORT_309_data = 32'h3f63c32a;
  assign cosLUT_MPORT_309_addr = 11'h135;
  assign cosLUT_MPORT_309_mask = 1'h1;
  assign cosLUT_MPORT_309_en = reset;
  assign cosLUT_MPORT_310_data = 32'h3f639530;
  assign cosLUT_MPORT_310_addr = 11'h136;
  assign cosLUT_MPORT_310_mask = 1'h1;
  assign cosLUT_MPORT_310_en = reset;
  assign cosLUT_MPORT_311_data = 32'h3f636713;
  assign cosLUT_MPORT_311_addr = 11'h137;
  assign cosLUT_MPORT_311_mask = 1'h1;
  assign cosLUT_MPORT_311_en = reset;
  assign cosLUT_MPORT_312_data = 32'h3f6338d3;
  assign cosLUT_MPORT_312_addr = 11'h138;
  assign cosLUT_MPORT_312_mask = 1'h1;
  assign cosLUT_MPORT_312_en = reset;
  assign cosLUT_MPORT_313_data = 32'h3f630a6f;
  assign cosLUT_MPORT_313_addr = 11'h139;
  assign cosLUT_MPORT_313_mask = 1'h1;
  assign cosLUT_MPORT_313_en = reset;
  assign cosLUT_MPORT_314_data = 32'h3f62dbe9;
  assign cosLUT_MPORT_314_addr = 11'h13a;
  assign cosLUT_MPORT_314_mask = 1'h1;
  assign cosLUT_MPORT_314_en = reset;
  assign cosLUT_MPORT_315_data = 32'h3f62ad3f;
  assign cosLUT_MPORT_315_addr = 11'h13b;
  assign cosLUT_MPORT_315_mask = 1'h1;
  assign cosLUT_MPORT_315_en = reset;
  assign cosLUT_MPORT_316_data = 32'h3f627e73;
  assign cosLUT_MPORT_316_addr = 11'h13c;
  assign cosLUT_MPORT_316_mask = 1'h1;
  assign cosLUT_MPORT_316_en = reset;
  assign cosLUT_MPORT_317_data = 32'h3f624f83;
  assign cosLUT_MPORT_317_addr = 11'h13d;
  assign cosLUT_MPORT_317_mask = 1'h1;
  assign cosLUT_MPORT_317_en = reset;
  assign cosLUT_MPORT_318_data = 32'h3f622071;
  assign cosLUT_MPORT_318_addr = 11'h13e;
  assign cosLUT_MPORT_318_mask = 1'h1;
  assign cosLUT_MPORT_318_en = reset;
  assign cosLUT_MPORT_319_data = 32'h3f61f13c;
  assign cosLUT_MPORT_319_addr = 11'h13f;
  assign cosLUT_MPORT_319_mask = 1'h1;
  assign cosLUT_MPORT_319_en = reset;
  assign cosLUT_MPORT_320_data = 32'h3f61c1e3;
  assign cosLUT_MPORT_320_addr = 11'h140;
  assign cosLUT_MPORT_320_mask = 1'h1;
  assign cosLUT_MPORT_320_en = reset;
  assign cosLUT_MPORT_321_data = 32'h3f619268;
  assign cosLUT_MPORT_321_addr = 11'h141;
  assign cosLUT_MPORT_321_mask = 1'h1;
  assign cosLUT_MPORT_321_en = reset;
  assign cosLUT_MPORT_322_data = 32'h3f6162cb;
  assign cosLUT_MPORT_322_addr = 11'h142;
  assign cosLUT_MPORT_322_mask = 1'h1;
  assign cosLUT_MPORT_322_en = reset;
  assign cosLUT_MPORT_323_data = 32'h3f61330a;
  assign cosLUT_MPORT_323_addr = 11'h143;
  assign cosLUT_MPORT_323_mask = 1'h1;
  assign cosLUT_MPORT_323_en = reset;
  assign cosLUT_MPORT_324_data = 32'h3f610327;
  assign cosLUT_MPORT_324_addr = 11'h144;
  assign cosLUT_MPORT_324_mask = 1'h1;
  assign cosLUT_MPORT_324_en = reset;
  assign cosLUT_MPORT_325_data = 32'h3f60d321;
  assign cosLUT_MPORT_325_addr = 11'h145;
  assign cosLUT_MPORT_325_mask = 1'h1;
  assign cosLUT_MPORT_325_en = reset;
  assign cosLUT_MPORT_326_data = 32'h3f60a2f8;
  assign cosLUT_MPORT_326_addr = 11'h146;
  assign cosLUT_MPORT_326_mask = 1'h1;
  assign cosLUT_MPORT_326_en = reset;
  assign cosLUT_MPORT_327_data = 32'h3f6072ad;
  assign cosLUT_MPORT_327_addr = 11'h147;
  assign cosLUT_MPORT_327_mask = 1'h1;
  assign cosLUT_MPORT_327_en = reset;
  assign cosLUT_MPORT_328_data = 32'h3f60423f;
  assign cosLUT_MPORT_328_addr = 11'h148;
  assign cosLUT_MPORT_328_mask = 1'h1;
  assign cosLUT_MPORT_328_en = reset;
  assign cosLUT_MPORT_329_data = 32'h3f6011af;
  assign cosLUT_MPORT_329_addr = 11'h149;
  assign cosLUT_MPORT_329_mask = 1'h1;
  assign cosLUT_MPORT_329_en = reset;
  assign cosLUT_MPORT_330_data = 32'h3f5fe0fb;
  assign cosLUT_MPORT_330_addr = 11'h14a;
  assign cosLUT_MPORT_330_mask = 1'h1;
  assign cosLUT_MPORT_330_en = reset;
  assign cosLUT_MPORT_331_data = 32'h3f5fb026;
  assign cosLUT_MPORT_331_addr = 11'h14b;
  assign cosLUT_MPORT_331_mask = 1'h1;
  assign cosLUT_MPORT_331_en = reset;
  assign cosLUT_MPORT_332_data = 32'h3f5f7f2e;
  assign cosLUT_MPORT_332_addr = 11'h14c;
  assign cosLUT_MPORT_332_mask = 1'h1;
  assign cosLUT_MPORT_332_en = reset;
  assign cosLUT_MPORT_333_data = 32'h3f5f4e13;
  assign cosLUT_MPORT_333_addr = 11'h14d;
  assign cosLUT_MPORT_333_mask = 1'h1;
  assign cosLUT_MPORT_333_en = reset;
  assign cosLUT_MPORT_334_data = 32'h3f5f1cd6;
  assign cosLUT_MPORT_334_addr = 11'h14e;
  assign cosLUT_MPORT_334_mask = 1'h1;
  assign cosLUT_MPORT_334_en = reset;
  assign cosLUT_MPORT_335_data = 32'h3f5eeb76;
  assign cosLUT_MPORT_335_addr = 11'h14f;
  assign cosLUT_MPORT_335_mask = 1'h1;
  assign cosLUT_MPORT_335_en = reset;
  assign cosLUT_MPORT_336_data = 32'h3f5eb9f4;
  assign cosLUT_MPORT_336_addr = 11'h150;
  assign cosLUT_MPORT_336_mask = 1'h1;
  assign cosLUT_MPORT_336_en = reset;
  assign cosLUT_MPORT_337_data = 32'h3f5e8850;
  assign cosLUT_MPORT_337_addr = 11'h151;
  assign cosLUT_MPORT_337_mask = 1'h1;
  assign cosLUT_MPORT_337_en = reset;
  assign cosLUT_MPORT_338_data = 32'h3f5e568a;
  assign cosLUT_MPORT_338_addr = 11'h152;
  assign cosLUT_MPORT_338_mask = 1'h1;
  assign cosLUT_MPORT_338_en = reset;
  assign cosLUT_MPORT_339_data = 32'h3f5e24a1;
  assign cosLUT_MPORT_339_addr = 11'h153;
  assign cosLUT_MPORT_339_mask = 1'h1;
  assign cosLUT_MPORT_339_en = reset;
  assign cosLUT_MPORT_340_data = 32'h3f5df295;
  assign cosLUT_MPORT_340_addr = 11'h154;
  assign cosLUT_MPORT_340_mask = 1'h1;
  assign cosLUT_MPORT_340_en = reset;
  assign cosLUT_MPORT_341_data = 32'h3f5dc068;
  assign cosLUT_MPORT_341_addr = 11'h155;
  assign cosLUT_MPORT_341_mask = 1'h1;
  assign cosLUT_MPORT_341_en = reset;
  assign cosLUT_MPORT_342_data = 32'h3f5d8e18;
  assign cosLUT_MPORT_342_addr = 11'h156;
  assign cosLUT_MPORT_342_mask = 1'h1;
  assign cosLUT_MPORT_342_en = reset;
  assign cosLUT_MPORT_343_data = 32'h3f5d5ba6;
  assign cosLUT_MPORT_343_addr = 11'h157;
  assign cosLUT_MPORT_343_mask = 1'h1;
  assign cosLUT_MPORT_343_en = reset;
  assign cosLUT_MPORT_344_data = 32'h3f5d2912;
  assign cosLUT_MPORT_344_addr = 11'h158;
  assign cosLUT_MPORT_344_mask = 1'h1;
  assign cosLUT_MPORT_344_en = reset;
  assign cosLUT_MPORT_345_data = 32'h3f5cf65c;
  assign cosLUT_MPORT_345_addr = 11'h159;
  assign cosLUT_MPORT_345_mask = 1'h1;
  assign cosLUT_MPORT_345_en = reset;
  assign cosLUT_MPORT_346_data = 32'h3f5cc384;
  assign cosLUT_MPORT_346_addr = 11'h15a;
  assign cosLUT_MPORT_346_mask = 1'h1;
  assign cosLUT_MPORT_346_en = reset;
  assign cosLUT_MPORT_347_data = 32'h3f5c908a;
  assign cosLUT_MPORT_347_addr = 11'h15b;
  assign cosLUT_MPORT_347_mask = 1'h1;
  assign cosLUT_MPORT_347_en = reset;
  assign cosLUT_MPORT_348_data = 32'h3f5c5d6e;
  assign cosLUT_MPORT_348_addr = 11'h15c;
  assign cosLUT_MPORT_348_mask = 1'h1;
  assign cosLUT_MPORT_348_en = reset;
  assign cosLUT_MPORT_349_data = 32'h3f5c2a2f;
  assign cosLUT_MPORT_349_addr = 11'h15d;
  assign cosLUT_MPORT_349_mask = 1'h1;
  assign cosLUT_MPORT_349_en = reset;
  assign cosLUT_MPORT_350_data = 32'h3f5bf6cf;
  assign cosLUT_MPORT_350_addr = 11'h15e;
  assign cosLUT_MPORT_350_mask = 1'h1;
  assign cosLUT_MPORT_350_en = reset;
  assign cosLUT_MPORT_351_data = 32'h3f5bc34d;
  assign cosLUT_MPORT_351_addr = 11'h15f;
  assign cosLUT_MPORT_351_mask = 1'h1;
  assign cosLUT_MPORT_351_en = reset;
  assign cosLUT_MPORT_352_data = 32'h3f5b8fa9;
  assign cosLUT_MPORT_352_addr = 11'h160;
  assign cosLUT_MPORT_352_mask = 1'h1;
  assign cosLUT_MPORT_352_en = reset;
  assign cosLUT_MPORT_353_data = 32'h3f5b5be3;
  assign cosLUT_MPORT_353_addr = 11'h161;
  assign cosLUT_MPORT_353_mask = 1'h1;
  assign cosLUT_MPORT_353_en = reset;
  assign cosLUT_MPORT_354_data = 32'h3f5b27fb;
  assign cosLUT_MPORT_354_addr = 11'h162;
  assign cosLUT_MPORT_354_mask = 1'h1;
  assign cosLUT_MPORT_354_en = reset;
  assign cosLUT_MPORT_355_data = 32'h3f5af3f1;
  assign cosLUT_MPORT_355_addr = 11'h163;
  assign cosLUT_MPORT_355_mask = 1'h1;
  assign cosLUT_MPORT_355_en = reset;
  assign cosLUT_MPORT_356_data = 32'h3f5abfc6;
  assign cosLUT_MPORT_356_addr = 11'h164;
  assign cosLUT_MPORT_356_mask = 1'h1;
  assign cosLUT_MPORT_356_en = reset;
  assign cosLUT_MPORT_357_data = 32'h3f5a8b79;
  assign cosLUT_MPORT_357_addr = 11'h165;
  assign cosLUT_MPORT_357_mask = 1'h1;
  assign cosLUT_MPORT_357_en = reset;
  assign cosLUT_MPORT_358_data = 32'h3f5a570a;
  assign cosLUT_MPORT_358_addr = 11'h166;
  assign cosLUT_MPORT_358_mask = 1'h1;
  assign cosLUT_MPORT_358_en = reset;
  assign cosLUT_MPORT_359_data = 32'h3f5a2279;
  assign cosLUT_MPORT_359_addr = 11'h167;
  assign cosLUT_MPORT_359_mask = 1'h1;
  assign cosLUT_MPORT_359_en = reset;
  assign cosLUT_MPORT_360_data = 32'h3f59edc7;
  assign cosLUT_MPORT_360_addr = 11'h168;
  assign cosLUT_MPORT_360_mask = 1'h1;
  assign cosLUT_MPORT_360_en = reset;
  assign cosLUT_MPORT_361_data = 32'h3f59b8f3;
  assign cosLUT_MPORT_361_addr = 11'h169;
  assign cosLUT_MPORT_361_mask = 1'h1;
  assign cosLUT_MPORT_361_en = reset;
  assign cosLUT_MPORT_362_data = 32'h3f5983fe;
  assign cosLUT_MPORT_362_addr = 11'h16a;
  assign cosLUT_MPORT_362_mask = 1'h1;
  assign cosLUT_MPORT_362_en = reset;
  assign cosLUT_MPORT_363_data = 32'h3f594ee7;
  assign cosLUT_MPORT_363_addr = 11'h16b;
  assign cosLUT_MPORT_363_mask = 1'h1;
  assign cosLUT_MPORT_363_en = reset;
  assign cosLUT_MPORT_364_data = 32'h3f5919ae;
  assign cosLUT_MPORT_364_addr = 11'h16c;
  assign cosLUT_MPORT_364_mask = 1'h1;
  assign cosLUT_MPORT_364_en = reset;
  assign cosLUT_MPORT_365_data = 32'h3f58e454;
  assign cosLUT_MPORT_365_addr = 11'h16d;
  assign cosLUT_MPORT_365_mask = 1'h1;
  assign cosLUT_MPORT_365_en = reset;
  assign cosLUT_MPORT_366_data = 32'h3f58aed9;
  assign cosLUT_MPORT_366_addr = 11'h16e;
  assign cosLUT_MPORT_366_mask = 1'h1;
  assign cosLUT_MPORT_366_en = reset;
  assign cosLUT_MPORT_367_data = 32'h3f58793c;
  assign cosLUT_MPORT_367_addr = 11'h16f;
  assign cosLUT_MPORT_367_mask = 1'h1;
  assign cosLUT_MPORT_367_en = reset;
  assign cosLUT_MPORT_368_data = 32'h3f58437d;
  assign cosLUT_MPORT_368_addr = 11'h170;
  assign cosLUT_MPORT_368_mask = 1'h1;
  assign cosLUT_MPORT_368_en = reset;
  assign cosLUT_MPORT_369_data = 32'h3f580d9e;
  assign cosLUT_MPORT_369_addr = 11'h171;
  assign cosLUT_MPORT_369_mask = 1'h1;
  assign cosLUT_MPORT_369_en = reset;
  assign cosLUT_MPORT_370_data = 32'h3f57d79d;
  assign cosLUT_MPORT_370_addr = 11'h172;
  assign cosLUT_MPORT_370_mask = 1'h1;
  assign cosLUT_MPORT_370_en = reset;
  assign cosLUT_MPORT_371_data = 32'h3f57a17a;
  assign cosLUT_MPORT_371_addr = 11'h173;
  assign cosLUT_MPORT_371_mask = 1'h1;
  assign cosLUT_MPORT_371_en = reset;
  assign cosLUT_MPORT_372_data = 32'h3f576b37;
  assign cosLUT_MPORT_372_addr = 11'h174;
  assign cosLUT_MPORT_372_mask = 1'h1;
  assign cosLUT_MPORT_372_en = reset;
  assign cosLUT_MPORT_373_data = 32'h3f5734d2;
  assign cosLUT_MPORT_373_addr = 11'h175;
  assign cosLUT_MPORT_373_mask = 1'h1;
  assign cosLUT_MPORT_373_en = reset;
  assign cosLUT_MPORT_374_data = 32'h3f56fe4c;
  assign cosLUT_MPORT_374_addr = 11'h176;
  assign cosLUT_MPORT_374_mask = 1'h1;
  assign cosLUT_MPORT_374_en = reset;
  assign cosLUT_MPORT_375_data = 32'h3f56c7a5;
  assign cosLUT_MPORT_375_addr = 11'h177;
  assign cosLUT_MPORT_375_mask = 1'h1;
  assign cosLUT_MPORT_375_en = reset;
  assign cosLUT_MPORT_376_data = 32'h3f5690dc;
  assign cosLUT_MPORT_376_addr = 11'h178;
  assign cosLUT_MPORT_376_mask = 1'h1;
  assign cosLUT_MPORT_376_en = reset;
  assign cosLUT_MPORT_377_data = 32'h3f5659f3;
  assign cosLUT_MPORT_377_addr = 11'h179;
  assign cosLUT_MPORT_377_mask = 1'h1;
  assign cosLUT_MPORT_377_en = reset;
  assign cosLUT_MPORT_378_data = 32'h3f5622e8;
  assign cosLUT_MPORT_378_addr = 11'h17a;
  assign cosLUT_MPORT_378_mask = 1'h1;
  assign cosLUT_MPORT_378_en = reset;
  assign cosLUT_MPORT_379_data = 32'h3f55ebbd;
  assign cosLUT_MPORT_379_addr = 11'h17b;
  assign cosLUT_MPORT_379_mask = 1'h1;
  assign cosLUT_MPORT_379_en = reset;
  assign cosLUT_MPORT_380_data = 32'h3f55b470;
  assign cosLUT_MPORT_380_addr = 11'h17c;
  assign cosLUT_MPORT_380_mask = 1'h1;
  assign cosLUT_MPORT_380_en = reset;
  assign cosLUT_MPORT_381_data = 32'h3f557d02;
  assign cosLUT_MPORT_381_addr = 11'h17d;
  assign cosLUT_MPORT_381_mask = 1'h1;
  assign cosLUT_MPORT_381_en = reset;
  assign cosLUT_MPORT_382_data = 32'h3f554574;
  assign cosLUT_MPORT_382_addr = 11'h17e;
  assign cosLUT_MPORT_382_mask = 1'h1;
  assign cosLUT_MPORT_382_en = reset;
  assign cosLUT_MPORT_383_data = 32'h3f550dc5;
  assign cosLUT_MPORT_383_addr = 11'h17f;
  assign cosLUT_MPORT_383_mask = 1'h1;
  assign cosLUT_MPORT_383_en = reset;
  assign cosLUT_MPORT_384_data = 32'h3f54d5f4;
  assign cosLUT_MPORT_384_addr = 11'h180;
  assign cosLUT_MPORT_384_mask = 1'h1;
  assign cosLUT_MPORT_384_en = reset;
  assign cosLUT_MPORT_385_data = 32'h3f549e03;
  assign cosLUT_MPORT_385_addr = 11'h181;
  assign cosLUT_MPORT_385_mask = 1'h1;
  assign cosLUT_MPORT_385_en = reset;
  assign cosLUT_MPORT_386_data = 32'h3f5465f1;
  assign cosLUT_MPORT_386_addr = 11'h182;
  assign cosLUT_MPORT_386_mask = 1'h1;
  assign cosLUT_MPORT_386_en = reset;
  assign cosLUT_MPORT_387_data = 32'h3f542dbf;
  assign cosLUT_MPORT_387_addr = 11'h183;
  assign cosLUT_MPORT_387_mask = 1'h1;
  assign cosLUT_MPORT_387_en = reset;
  assign cosLUT_MPORT_388_data = 32'h3f53f56b;
  assign cosLUT_MPORT_388_addr = 11'h184;
  assign cosLUT_MPORT_388_mask = 1'h1;
  assign cosLUT_MPORT_388_en = reset;
  assign cosLUT_MPORT_389_data = 32'h3f53bcf7;
  assign cosLUT_MPORT_389_addr = 11'h185;
  assign cosLUT_MPORT_389_mask = 1'h1;
  assign cosLUT_MPORT_389_en = reset;
  assign cosLUT_MPORT_390_data = 32'h3f538462;
  assign cosLUT_MPORT_390_addr = 11'h186;
  assign cosLUT_MPORT_390_mask = 1'h1;
  assign cosLUT_MPORT_390_en = reset;
  assign cosLUT_MPORT_391_data = 32'h3f534bad;
  assign cosLUT_MPORT_391_addr = 11'h187;
  assign cosLUT_MPORT_391_mask = 1'h1;
  assign cosLUT_MPORT_391_en = reset;
  assign cosLUT_MPORT_392_data = 32'h3f5312d7;
  assign cosLUT_MPORT_392_addr = 11'h188;
  assign cosLUT_MPORT_392_mask = 1'h1;
  assign cosLUT_MPORT_392_en = reset;
  assign cosLUT_MPORT_393_data = 32'h3f52d9e0;
  assign cosLUT_MPORT_393_addr = 11'h189;
  assign cosLUT_MPORT_393_mask = 1'h1;
  assign cosLUT_MPORT_393_en = reset;
  assign cosLUT_MPORT_394_data = 32'h3f52a0c9;
  assign cosLUT_MPORT_394_addr = 11'h18a;
  assign cosLUT_MPORT_394_mask = 1'h1;
  assign cosLUT_MPORT_394_en = reset;
  assign cosLUT_MPORT_395_data = 32'h3f526792;
  assign cosLUT_MPORT_395_addr = 11'h18b;
  assign cosLUT_MPORT_395_mask = 1'h1;
  assign cosLUT_MPORT_395_en = reset;
  assign cosLUT_MPORT_396_data = 32'h3f522e3a;
  assign cosLUT_MPORT_396_addr = 11'h18c;
  assign cosLUT_MPORT_396_mask = 1'h1;
  assign cosLUT_MPORT_396_en = reset;
  assign cosLUT_MPORT_397_data = 32'h3f51f4c1;
  assign cosLUT_MPORT_397_addr = 11'h18d;
  assign cosLUT_MPORT_397_mask = 1'h1;
  assign cosLUT_MPORT_397_en = reset;
  assign cosLUT_MPORT_398_data = 32'h3f51bb28;
  assign cosLUT_MPORT_398_addr = 11'h18e;
  assign cosLUT_MPORT_398_mask = 1'h1;
  assign cosLUT_MPORT_398_en = reset;
  assign cosLUT_MPORT_399_data = 32'h3f51816f;
  assign cosLUT_MPORT_399_addr = 11'h18f;
  assign cosLUT_MPORT_399_mask = 1'h1;
  assign cosLUT_MPORT_399_en = reset;
  assign cosLUT_MPORT_400_data = 32'h3f514795;
  assign cosLUT_MPORT_400_addr = 11'h190;
  assign cosLUT_MPORT_400_mask = 1'h1;
  assign cosLUT_MPORT_400_en = reset;
  assign cosLUT_MPORT_401_data = 32'h3f510d9b;
  assign cosLUT_MPORT_401_addr = 11'h191;
  assign cosLUT_MPORT_401_mask = 1'h1;
  assign cosLUT_MPORT_401_en = reset;
  assign cosLUT_MPORT_402_data = 32'h3f50d381;
  assign cosLUT_MPORT_402_addr = 11'h192;
  assign cosLUT_MPORT_402_mask = 1'h1;
  assign cosLUT_MPORT_402_en = reset;
  assign cosLUT_MPORT_403_data = 32'h3f509947;
  assign cosLUT_MPORT_403_addr = 11'h193;
  assign cosLUT_MPORT_403_mask = 1'h1;
  assign cosLUT_MPORT_403_en = reset;
  assign cosLUT_MPORT_404_data = 32'h3f505eec;
  assign cosLUT_MPORT_404_addr = 11'h194;
  assign cosLUT_MPORT_404_mask = 1'h1;
  assign cosLUT_MPORT_404_en = reset;
  assign cosLUT_MPORT_405_data = 32'h3f502472;
  assign cosLUT_MPORT_405_addr = 11'h195;
  assign cosLUT_MPORT_405_mask = 1'h1;
  assign cosLUT_MPORT_405_en = reset;
  assign cosLUT_MPORT_406_data = 32'h3f4fe9d7;
  assign cosLUT_MPORT_406_addr = 11'h196;
  assign cosLUT_MPORT_406_mask = 1'h1;
  assign cosLUT_MPORT_406_en = reset;
  assign cosLUT_MPORT_407_data = 32'h3f4faf1c;
  assign cosLUT_MPORT_407_addr = 11'h197;
  assign cosLUT_MPORT_407_mask = 1'h1;
  assign cosLUT_MPORT_407_en = reset;
  assign cosLUT_MPORT_408_data = 32'h3f4f7441;
  assign cosLUT_MPORT_408_addr = 11'h198;
  assign cosLUT_MPORT_408_mask = 1'h1;
  assign cosLUT_MPORT_408_en = reset;
  assign cosLUT_MPORT_409_data = 32'h3f4f3946;
  assign cosLUT_MPORT_409_addr = 11'h199;
  assign cosLUT_MPORT_409_mask = 1'h1;
  assign cosLUT_MPORT_409_en = reset;
  assign cosLUT_MPORT_410_data = 32'h3f4efe2b;
  assign cosLUT_MPORT_410_addr = 11'h19a;
  assign cosLUT_MPORT_410_mask = 1'h1;
  assign cosLUT_MPORT_410_en = reset;
  assign cosLUT_MPORT_411_data = 32'h3f4ec2f1;
  assign cosLUT_MPORT_411_addr = 11'h19b;
  assign cosLUT_MPORT_411_mask = 1'h1;
  assign cosLUT_MPORT_411_en = reset;
  assign cosLUT_MPORT_412_data = 32'h3f4e8796;
  assign cosLUT_MPORT_412_addr = 11'h19c;
  assign cosLUT_MPORT_412_mask = 1'h1;
  assign cosLUT_MPORT_412_en = reset;
  assign cosLUT_MPORT_413_data = 32'h3f4e4c1b;
  assign cosLUT_MPORT_413_addr = 11'h19d;
  assign cosLUT_MPORT_413_mask = 1'h1;
  assign cosLUT_MPORT_413_en = reset;
  assign cosLUT_MPORT_414_data = 32'h3f4e1081;
  assign cosLUT_MPORT_414_addr = 11'h19e;
  assign cosLUT_MPORT_414_mask = 1'h1;
  assign cosLUT_MPORT_414_en = reset;
  assign cosLUT_MPORT_415_data = 32'h3f4dd4c7;
  assign cosLUT_MPORT_415_addr = 11'h19f;
  assign cosLUT_MPORT_415_mask = 1'h1;
  assign cosLUT_MPORT_415_en = reset;
  assign cosLUT_MPORT_416_data = 32'h3f4d98ed;
  assign cosLUT_MPORT_416_addr = 11'h1a0;
  assign cosLUT_MPORT_416_mask = 1'h1;
  assign cosLUT_MPORT_416_en = reset;
  assign cosLUT_MPORT_417_data = 32'h3f4d5cf3;
  assign cosLUT_MPORT_417_addr = 11'h1a1;
  assign cosLUT_MPORT_417_mask = 1'h1;
  assign cosLUT_MPORT_417_en = reset;
  assign cosLUT_MPORT_418_data = 32'h3f4d20da;
  assign cosLUT_MPORT_418_addr = 11'h1a2;
  assign cosLUT_MPORT_418_mask = 1'h1;
  assign cosLUT_MPORT_418_en = reset;
  assign cosLUT_MPORT_419_data = 32'h3f4ce4a1;
  assign cosLUT_MPORT_419_addr = 11'h1a3;
  assign cosLUT_MPORT_419_mask = 1'h1;
  assign cosLUT_MPORT_419_en = reset;
  assign cosLUT_MPORT_420_data = 32'h3f4ca848;
  assign cosLUT_MPORT_420_addr = 11'h1a4;
  assign cosLUT_MPORT_420_mask = 1'h1;
  assign cosLUT_MPORT_420_en = reset;
  assign cosLUT_MPORT_421_data = 32'h3f4c6bd0;
  assign cosLUT_MPORT_421_addr = 11'h1a5;
  assign cosLUT_MPORT_421_mask = 1'h1;
  assign cosLUT_MPORT_421_en = reset;
  assign cosLUT_MPORT_422_data = 32'h3f4c2f38;
  assign cosLUT_MPORT_422_addr = 11'h1a6;
  assign cosLUT_MPORT_422_mask = 1'h1;
  assign cosLUT_MPORT_422_en = reset;
  assign cosLUT_MPORT_423_data = 32'h3f4bf281;
  assign cosLUT_MPORT_423_addr = 11'h1a7;
  assign cosLUT_MPORT_423_mask = 1'h1;
  assign cosLUT_MPORT_423_en = reset;
  assign cosLUT_MPORT_424_data = 32'h3f4bb5aa;
  assign cosLUT_MPORT_424_addr = 11'h1a8;
  assign cosLUT_MPORT_424_mask = 1'h1;
  assign cosLUT_MPORT_424_en = reset;
  assign cosLUT_MPORT_425_data = 32'h3f4b78b4;
  assign cosLUT_MPORT_425_addr = 11'h1a9;
  assign cosLUT_MPORT_425_mask = 1'h1;
  assign cosLUT_MPORT_425_en = reset;
  assign cosLUT_MPORT_426_data = 32'h3f4b3b9e;
  assign cosLUT_MPORT_426_addr = 11'h1aa;
  assign cosLUT_MPORT_426_mask = 1'h1;
  assign cosLUT_MPORT_426_en = reset;
  assign cosLUT_MPORT_427_data = 32'h3f4afe69;
  assign cosLUT_MPORT_427_addr = 11'h1ab;
  assign cosLUT_MPORT_427_mask = 1'h1;
  assign cosLUT_MPORT_427_en = reset;
  assign cosLUT_MPORT_428_data = 32'h3f4ac115;
  assign cosLUT_MPORT_428_addr = 11'h1ac;
  assign cosLUT_MPORT_428_mask = 1'h1;
  assign cosLUT_MPORT_428_en = reset;
  assign cosLUT_MPORT_429_data = 32'h3f4a83a2;
  assign cosLUT_MPORT_429_addr = 11'h1ad;
  assign cosLUT_MPORT_429_mask = 1'h1;
  assign cosLUT_MPORT_429_en = reset;
  assign cosLUT_MPORT_430_data = 32'h3f4a460f;
  assign cosLUT_MPORT_430_addr = 11'h1ae;
  assign cosLUT_MPORT_430_mask = 1'h1;
  assign cosLUT_MPORT_430_en = reset;
  assign cosLUT_MPORT_431_data = 32'h3f4a085d;
  assign cosLUT_MPORT_431_addr = 11'h1af;
  assign cosLUT_MPORT_431_mask = 1'h1;
  assign cosLUT_MPORT_431_en = reset;
  assign cosLUT_MPORT_432_data = 32'h3f49ca8c;
  assign cosLUT_MPORT_432_addr = 11'h1b0;
  assign cosLUT_MPORT_432_mask = 1'h1;
  assign cosLUT_MPORT_432_en = reset;
  assign cosLUT_MPORT_433_data = 32'h3f498c9c;
  assign cosLUT_MPORT_433_addr = 11'h1b1;
  assign cosLUT_MPORT_433_mask = 1'h1;
  assign cosLUT_MPORT_433_en = reset;
  assign cosLUT_MPORT_434_data = 32'h3f494e8c;
  assign cosLUT_MPORT_434_addr = 11'h1b2;
  assign cosLUT_MPORT_434_mask = 1'h1;
  assign cosLUT_MPORT_434_en = reset;
  assign cosLUT_MPORT_435_data = 32'h3f49105e;
  assign cosLUT_MPORT_435_addr = 11'h1b3;
  assign cosLUT_MPORT_435_mask = 1'h1;
  assign cosLUT_MPORT_435_en = reset;
  assign cosLUT_MPORT_436_data = 32'h3f48d210;
  assign cosLUT_MPORT_436_addr = 11'h1b4;
  assign cosLUT_MPORT_436_mask = 1'h1;
  assign cosLUT_MPORT_436_en = reset;
  assign cosLUT_MPORT_437_data = 32'h3f4893a4;
  assign cosLUT_MPORT_437_addr = 11'h1b5;
  assign cosLUT_MPORT_437_mask = 1'h1;
  assign cosLUT_MPORT_437_en = reset;
  assign cosLUT_MPORT_438_data = 32'h3f485518;
  assign cosLUT_MPORT_438_addr = 11'h1b6;
  assign cosLUT_MPORT_438_mask = 1'h1;
  assign cosLUT_MPORT_438_en = reset;
  assign cosLUT_MPORT_439_data = 32'h3f48166e;
  assign cosLUT_MPORT_439_addr = 11'h1b7;
  assign cosLUT_MPORT_439_mask = 1'h1;
  assign cosLUT_MPORT_439_en = reset;
  assign cosLUT_MPORT_440_data = 32'h3f47d7a5;
  assign cosLUT_MPORT_440_addr = 11'h1b8;
  assign cosLUT_MPORT_440_mask = 1'h1;
  assign cosLUT_MPORT_440_en = reset;
  assign cosLUT_MPORT_441_data = 32'h3f4798bd;
  assign cosLUT_MPORT_441_addr = 11'h1b9;
  assign cosLUT_MPORT_441_mask = 1'h1;
  assign cosLUT_MPORT_441_en = reset;
  assign cosLUT_MPORT_442_data = 32'h3f4759b6;
  assign cosLUT_MPORT_442_addr = 11'h1ba;
  assign cosLUT_MPORT_442_mask = 1'h1;
  assign cosLUT_MPORT_442_en = reset;
  assign cosLUT_MPORT_443_data = 32'h3f471a91;
  assign cosLUT_MPORT_443_addr = 11'h1bb;
  assign cosLUT_MPORT_443_mask = 1'h1;
  assign cosLUT_MPORT_443_en = reset;
  assign cosLUT_MPORT_444_data = 32'h3f46db4c;
  assign cosLUT_MPORT_444_addr = 11'h1bc;
  assign cosLUT_MPORT_444_mask = 1'h1;
  assign cosLUT_MPORT_444_en = reset;
  assign cosLUT_MPORT_445_data = 32'h3f469bea;
  assign cosLUT_MPORT_445_addr = 11'h1bd;
  assign cosLUT_MPORT_445_mask = 1'h1;
  assign cosLUT_MPORT_445_en = reset;
  assign cosLUT_MPORT_446_data = 32'h3f465c68;
  assign cosLUT_MPORT_446_addr = 11'h1be;
  assign cosLUT_MPORT_446_mask = 1'h1;
  assign cosLUT_MPORT_446_en = reset;
  assign cosLUT_MPORT_447_data = 32'h3f461cc8;
  assign cosLUT_MPORT_447_addr = 11'h1bf;
  assign cosLUT_MPORT_447_mask = 1'h1;
  assign cosLUT_MPORT_447_en = reset;
  assign cosLUT_MPORT_448_data = 32'h3f45dd09;
  assign cosLUT_MPORT_448_addr = 11'h1c0;
  assign cosLUT_MPORT_448_mask = 1'h1;
  assign cosLUT_MPORT_448_en = reset;
  assign cosLUT_MPORT_449_data = 32'h3f459d2c;
  assign cosLUT_MPORT_449_addr = 11'h1c1;
  assign cosLUT_MPORT_449_mask = 1'h1;
  assign cosLUT_MPORT_449_en = reset;
  assign cosLUT_MPORT_450_data = 32'h3f455d30;
  assign cosLUT_MPORT_450_addr = 11'h1c2;
  assign cosLUT_MPORT_450_mask = 1'h1;
  assign cosLUT_MPORT_450_en = reset;
  assign cosLUT_MPORT_451_data = 32'h3f451d16;
  assign cosLUT_MPORT_451_addr = 11'h1c3;
  assign cosLUT_MPORT_451_mask = 1'h1;
  assign cosLUT_MPORT_451_en = reset;
  assign cosLUT_MPORT_452_data = 32'h3f44dcdd;
  assign cosLUT_MPORT_452_addr = 11'h1c4;
  assign cosLUT_MPORT_452_mask = 1'h1;
  assign cosLUT_MPORT_452_en = reset;
  assign cosLUT_MPORT_453_data = 32'h3f449c86;
  assign cosLUT_MPORT_453_addr = 11'h1c5;
  assign cosLUT_MPORT_453_mask = 1'h1;
  assign cosLUT_MPORT_453_en = reset;
  assign cosLUT_MPORT_454_data = 32'h3f445c11;
  assign cosLUT_MPORT_454_addr = 11'h1c6;
  assign cosLUT_MPORT_454_mask = 1'h1;
  assign cosLUT_MPORT_454_en = reset;
  assign cosLUT_MPORT_455_data = 32'h3f441b7d;
  assign cosLUT_MPORT_455_addr = 11'h1c7;
  assign cosLUT_MPORT_455_mask = 1'h1;
  assign cosLUT_MPORT_455_en = reset;
  assign cosLUT_MPORT_456_data = 32'h3f43dacb;
  assign cosLUT_MPORT_456_addr = 11'h1c8;
  assign cosLUT_MPORT_456_mask = 1'h1;
  assign cosLUT_MPORT_456_en = reset;
  assign cosLUT_MPORT_457_data = 32'h3f4399fb;
  assign cosLUT_MPORT_457_addr = 11'h1c9;
  assign cosLUT_MPORT_457_mask = 1'h1;
  assign cosLUT_MPORT_457_en = reset;
  assign cosLUT_MPORT_458_data = 32'h3f43590d;
  assign cosLUT_MPORT_458_addr = 11'h1ca;
  assign cosLUT_MPORT_458_mask = 1'h1;
  assign cosLUT_MPORT_458_en = reset;
  assign cosLUT_MPORT_459_data = 32'h3f431800;
  assign cosLUT_MPORT_459_addr = 11'h1cb;
  assign cosLUT_MPORT_459_mask = 1'h1;
  assign cosLUT_MPORT_459_en = reset;
  assign cosLUT_MPORT_460_data = 32'h3f42d6d6;
  assign cosLUT_MPORT_460_addr = 11'h1cc;
  assign cosLUT_MPORT_460_mask = 1'h1;
  assign cosLUT_MPORT_460_en = reset;
  assign cosLUT_MPORT_461_data = 32'h3f42958d;
  assign cosLUT_MPORT_461_addr = 11'h1cd;
  assign cosLUT_MPORT_461_mask = 1'h1;
  assign cosLUT_MPORT_461_en = reset;
  assign cosLUT_MPORT_462_data = 32'h3f425427;
  assign cosLUT_MPORT_462_addr = 11'h1ce;
  assign cosLUT_MPORT_462_mask = 1'h1;
  assign cosLUT_MPORT_462_en = reset;
  assign cosLUT_MPORT_463_data = 32'h3f4212a2;
  assign cosLUT_MPORT_463_addr = 11'h1cf;
  assign cosLUT_MPORT_463_mask = 1'h1;
  assign cosLUT_MPORT_463_en = reset;
  assign cosLUT_MPORT_464_data = 32'h3f41d0ff;
  assign cosLUT_MPORT_464_addr = 11'h1d0;
  assign cosLUT_MPORT_464_mask = 1'h1;
  assign cosLUT_MPORT_464_en = reset;
  assign cosLUT_MPORT_465_data = 32'h3f418f3f;
  assign cosLUT_MPORT_465_addr = 11'h1d1;
  assign cosLUT_MPORT_465_mask = 1'h1;
  assign cosLUT_MPORT_465_en = reset;
  assign cosLUT_MPORT_466_data = 32'h3f414d61;
  assign cosLUT_MPORT_466_addr = 11'h1d2;
  assign cosLUT_MPORT_466_mask = 1'h1;
  assign cosLUT_MPORT_466_en = reset;
  assign cosLUT_MPORT_467_data = 32'h3f410b65;
  assign cosLUT_MPORT_467_addr = 11'h1d3;
  assign cosLUT_MPORT_467_mask = 1'h1;
  assign cosLUT_MPORT_467_en = reset;
  assign cosLUT_MPORT_468_data = 32'h3f40c94b;
  assign cosLUT_MPORT_468_addr = 11'h1d4;
  assign cosLUT_MPORT_468_mask = 1'h1;
  assign cosLUT_MPORT_468_en = reset;
  assign cosLUT_MPORT_469_data = 32'h3f408713;
  assign cosLUT_MPORT_469_addr = 11'h1d5;
  assign cosLUT_MPORT_469_mask = 1'h1;
  assign cosLUT_MPORT_469_en = reset;
  assign cosLUT_MPORT_470_data = 32'h3f4044be;
  assign cosLUT_MPORT_470_addr = 11'h1d6;
  assign cosLUT_MPORT_470_mask = 1'h1;
  assign cosLUT_MPORT_470_en = reset;
  assign cosLUT_MPORT_471_data = 32'h3f40024b;
  assign cosLUT_MPORT_471_addr = 11'h1d7;
  assign cosLUT_MPORT_471_mask = 1'h1;
  assign cosLUT_MPORT_471_en = reset;
  assign cosLUT_MPORT_472_data = 32'h3f3fbfba;
  assign cosLUT_MPORT_472_addr = 11'h1d8;
  assign cosLUT_MPORT_472_mask = 1'h1;
  assign cosLUT_MPORT_472_en = reset;
  assign cosLUT_MPORT_473_data = 32'h3f3f7d0c;
  assign cosLUT_MPORT_473_addr = 11'h1d9;
  assign cosLUT_MPORT_473_mask = 1'h1;
  assign cosLUT_MPORT_473_en = reset;
  assign cosLUT_MPORT_474_data = 32'h3f3f3a40;
  assign cosLUT_MPORT_474_addr = 11'h1da;
  assign cosLUT_MPORT_474_mask = 1'h1;
  assign cosLUT_MPORT_474_en = reset;
  assign cosLUT_MPORT_475_data = 32'h3f3ef757;
  assign cosLUT_MPORT_475_addr = 11'h1db;
  assign cosLUT_MPORT_475_mask = 1'h1;
  assign cosLUT_MPORT_475_en = reset;
  assign cosLUT_MPORT_476_data = 32'h3f3eb450;
  assign cosLUT_MPORT_476_addr = 11'h1dc;
  assign cosLUT_MPORT_476_mask = 1'h1;
  assign cosLUT_MPORT_476_en = reset;
  assign cosLUT_MPORT_477_data = 32'h3f3e712c;
  assign cosLUT_MPORT_477_addr = 11'h1dd;
  assign cosLUT_MPORT_477_mask = 1'h1;
  assign cosLUT_MPORT_477_en = reset;
  assign cosLUT_MPORT_478_data = 32'h3f3e2dea;
  assign cosLUT_MPORT_478_addr = 11'h1de;
  assign cosLUT_MPORT_478_mask = 1'h1;
  assign cosLUT_MPORT_478_en = reset;
  assign cosLUT_MPORT_479_data = 32'h3f3dea8b;
  assign cosLUT_MPORT_479_addr = 11'h1df;
  assign cosLUT_MPORT_479_mask = 1'h1;
  assign cosLUT_MPORT_479_en = reset;
  assign cosLUT_MPORT_480_data = 32'h3f3da70f;
  assign cosLUT_MPORT_480_addr = 11'h1e0;
  assign cosLUT_MPORT_480_mask = 1'h1;
  assign cosLUT_MPORT_480_en = reset;
  assign cosLUT_MPORT_481_data = 32'h3f3d6376;
  assign cosLUT_MPORT_481_addr = 11'h1e1;
  assign cosLUT_MPORT_481_mask = 1'h1;
  assign cosLUT_MPORT_481_en = reset;
  assign cosLUT_MPORT_482_data = 32'h3f3d1fbf;
  assign cosLUT_MPORT_482_addr = 11'h1e2;
  assign cosLUT_MPORT_482_mask = 1'h1;
  assign cosLUT_MPORT_482_en = reset;
  assign cosLUT_MPORT_483_data = 32'h3f3cdbeb;
  assign cosLUT_MPORT_483_addr = 11'h1e3;
  assign cosLUT_MPORT_483_mask = 1'h1;
  assign cosLUT_MPORT_483_en = reset;
  assign cosLUT_MPORT_484_data = 32'h3f3c97fa;
  assign cosLUT_MPORT_484_addr = 11'h1e4;
  assign cosLUT_MPORT_484_mask = 1'h1;
  assign cosLUT_MPORT_484_en = reset;
  assign cosLUT_MPORT_485_data = 32'h3f3c53ec;
  assign cosLUT_MPORT_485_addr = 11'h1e5;
  assign cosLUT_MPORT_485_mask = 1'h1;
  assign cosLUT_MPORT_485_en = reset;
  assign cosLUT_MPORT_486_data = 32'h3f3c0fc1;
  assign cosLUT_MPORT_486_addr = 11'h1e6;
  assign cosLUT_MPORT_486_mask = 1'h1;
  assign cosLUT_MPORT_486_en = reset;
  assign cosLUT_MPORT_487_data = 32'h3f3bcb79;
  assign cosLUT_MPORT_487_addr = 11'h1e7;
  assign cosLUT_MPORT_487_mask = 1'h1;
  assign cosLUT_MPORT_487_en = reset;
  assign cosLUT_MPORT_488_data = 32'h3f3b8713;
  assign cosLUT_MPORT_488_addr = 11'h1e8;
  assign cosLUT_MPORT_488_mask = 1'h1;
  assign cosLUT_MPORT_488_en = reset;
  assign cosLUT_MPORT_489_data = 32'h3f3b4291;
  assign cosLUT_MPORT_489_addr = 11'h1e9;
  assign cosLUT_MPORT_489_mask = 1'h1;
  assign cosLUT_MPORT_489_en = reset;
  assign cosLUT_MPORT_490_data = 32'h3f3afdf2;
  assign cosLUT_MPORT_490_addr = 11'h1ea;
  assign cosLUT_MPORT_490_mask = 1'h1;
  assign cosLUT_MPORT_490_en = reset;
  assign cosLUT_MPORT_491_data = 32'h3f3ab937;
  assign cosLUT_MPORT_491_addr = 11'h1eb;
  assign cosLUT_MPORT_491_mask = 1'h1;
  assign cosLUT_MPORT_491_en = reset;
  assign cosLUT_MPORT_492_data = 32'h3f3a745e;
  assign cosLUT_MPORT_492_addr = 11'h1ec;
  assign cosLUT_MPORT_492_mask = 1'h1;
  assign cosLUT_MPORT_492_en = reset;
  assign cosLUT_MPORT_493_data = 32'h3f3a2f68;
  assign cosLUT_MPORT_493_addr = 11'h1ed;
  assign cosLUT_MPORT_493_mask = 1'h1;
  assign cosLUT_MPORT_493_en = reset;
  assign cosLUT_MPORT_494_data = 32'h3f39ea56;
  assign cosLUT_MPORT_494_addr = 11'h1ee;
  assign cosLUT_MPORT_494_mask = 1'h1;
  assign cosLUT_MPORT_494_en = reset;
  assign cosLUT_MPORT_495_data = 32'h3f39a528;
  assign cosLUT_MPORT_495_addr = 11'h1ef;
  assign cosLUT_MPORT_495_mask = 1'h1;
  assign cosLUT_MPORT_495_en = reset;
  assign cosLUT_MPORT_496_data = 32'h3f395fdc;
  assign cosLUT_MPORT_496_addr = 11'h1f0;
  assign cosLUT_MPORT_496_mask = 1'h1;
  assign cosLUT_MPORT_496_en = reset;
  assign cosLUT_MPORT_497_data = 32'h3f391a74;
  assign cosLUT_MPORT_497_addr = 11'h1f1;
  assign cosLUT_MPORT_497_mask = 1'h1;
  assign cosLUT_MPORT_497_en = reset;
  assign cosLUT_MPORT_498_data = 32'h3f38d4ef;
  assign cosLUT_MPORT_498_addr = 11'h1f2;
  assign cosLUT_MPORT_498_mask = 1'h1;
  assign cosLUT_MPORT_498_en = reset;
  assign cosLUT_MPORT_499_data = 32'h3f388f4e;
  assign cosLUT_MPORT_499_addr = 11'h1f3;
  assign cosLUT_MPORT_499_mask = 1'h1;
  assign cosLUT_MPORT_499_en = reset;
  assign cosLUT_MPORT_500_data = 32'h3f384991;
  assign cosLUT_MPORT_500_addr = 11'h1f4;
  assign cosLUT_MPORT_500_mask = 1'h1;
  assign cosLUT_MPORT_500_en = reset;
  assign cosLUT_MPORT_501_data = 32'h3f3803b7;
  assign cosLUT_MPORT_501_addr = 11'h1f5;
  assign cosLUT_MPORT_501_mask = 1'h1;
  assign cosLUT_MPORT_501_en = reset;
  assign cosLUT_MPORT_502_data = 32'h3f37bdc0;
  assign cosLUT_MPORT_502_addr = 11'h1f6;
  assign cosLUT_MPORT_502_mask = 1'h1;
  assign cosLUT_MPORT_502_en = reset;
  assign cosLUT_MPORT_503_data = 32'h3f3777ad;
  assign cosLUT_MPORT_503_addr = 11'h1f7;
  assign cosLUT_MPORT_503_mask = 1'h1;
  assign cosLUT_MPORT_503_en = reset;
  assign cosLUT_MPORT_504_data = 32'h3f37317e;
  assign cosLUT_MPORT_504_addr = 11'h1f8;
  assign cosLUT_MPORT_504_mask = 1'h1;
  assign cosLUT_MPORT_504_en = reset;
  assign cosLUT_MPORT_505_data = 32'h3f36eb33;
  assign cosLUT_MPORT_505_addr = 11'h1f9;
  assign cosLUT_MPORT_505_mask = 1'h1;
  assign cosLUT_MPORT_505_en = reset;
  assign cosLUT_MPORT_506_data = 32'h3f36a4cb;
  assign cosLUT_MPORT_506_addr = 11'h1fa;
  assign cosLUT_MPORT_506_mask = 1'h1;
  assign cosLUT_MPORT_506_en = reset;
  assign cosLUT_MPORT_507_data = 32'h3f365e48;
  assign cosLUT_MPORT_507_addr = 11'h1fb;
  assign cosLUT_MPORT_507_mask = 1'h1;
  assign cosLUT_MPORT_507_en = reset;
  assign cosLUT_MPORT_508_data = 32'h3f3617a8;
  assign cosLUT_MPORT_508_addr = 11'h1fc;
  assign cosLUT_MPORT_508_mask = 1'h1;
  assign cosLUT_MPORT_508_en = reset;
  assign cosLUT_MPORT_509_data = 32'h3f35d0ec;
  assign cosLUT_MPORT_509_addr = 11'h1fd;
  assign cosLUT_MPORT_509_mask = 1'h1;
  assign cosLUT_MPORT_509_en = reset;
  assign cosLUT_MPORT_510_data = 32'h3f358a14;
  assign cosLUT_MPORT_510_addr = 11'h1fe;
  assign cosLUT_MPORT_510_mask = 1'h1;
  assign cosLUT_MPORT_510_en = reset;
  assign cosLUT_MPORT_511_data = 32'h3f354320;
  assign cosLUT_MPORT_511_addr = 11'h1ff;
  assign cosLUT_MPORT_511_mask = 1'h1;
  assign cosLUT_MPORT_511_en = reset;
  assign cosLUT_MPORT_512_data = 32'h3f34fc10;
  assign cosLUT_MPORT_512_addr = 11'h200;
  assign cosLUT_MPORT_512_mask = 1'h1;
  assign cosLUT_MPORT_512_en = reset;
  assign cosLUT_MPORT_513_data = 32'h3f34b4e4;
  assign cosLUT_MPORT_513_addr = 11'h201;
  assign cosLUT_MPORT_513_mask = 1'h1;
  assign cosLUT_MPORT_513_en = reset;
  assign cosLUT_MPORT_514_data = 32'h3f346d9c;
  assign cosLUT_MPORT_514_addr = 11'h202;
  assign cosLUT_MPORT_514_mask = 1'h1;
  assign cosLUT_MPORT_514_en = reset;
  assign cosLUT_MPORT_515_data = 32'h3f342638;
  assign cosLUT_MPORT_515_addr = 11'h203;
  assign cosLUT_MPORT_515_mask = 1'h1;
  assign cosLUT_MPORT_515_en = reset;
  assign cosLUT_MPORT_516_data = 32'h3f33deb9;
  assign cosLUT_MPORT_516_addr = 11'h204;
  assign cosLUT_MPORT_516_mask = 1'h1;
  assign cosLUT_MPORT_516_en = reset;
  assign cosLUT_MPORT_517_data = 32'h3f33971e;
  assign cosLUT_MPORT_517_addr = 11'h205;
  assign cosLUT_MPORT_517_mask = 1'h1;
  assign cosLUT_MPORT_517_en = reset;
  assign cosLUT_MPORT_518_data = 32'h3f334f67;
  assign cosLUT_MPORT_518_addr = 11'h206;
  assign cosLUT_MPORT_518_mask = 1'h1;
  assign cosLUT_MPORT_518_en = reset;
  assign cosLUT_MPORT_519_data = 32'h3f330794;
  assign cosLUT_MPORT_519_addr = 11'h207;
  assign cosLUT_MPORT_519_mask = 1'h1;
  assign cosLUT_MPORT_519_en = reset;
  assign cosLUT_MPORT_520_data = 32'h3f32bfa6;
  assign cosLUT_MPORT_520_addr = 11'h208;
  assign cosLUT_MPORT_520_mask = 1'h1;
  assign cosLUT_MPORT_520_en = reset;
  assign cosLUT_MPORT_521_data = 32'h3f32779c;
  assign cosLUT_MPORT_521_addr = 11'h209;
  assign cosLUT_MPORT_521_mask = 1'h1;
  assign cosLUT_MPORT_521_en = reset;
  assign cosLUT_MPORT_522_data = 32'h3f322f77;
  assign cosLUT_MPORT_522_addr = 11'h20a;
  assign cosLUT_MPORT_522_mask = 1'h1;
  assign cosLUT_MPORT_522_en = reset;
  assign cosLUT_MPORT_523_data = 32'h3f31e736;
  assign cosLUT_MPORT_523_addr = 11'h20b;
  assign cosLUT_MPORT_523_mask = 1'h1;
  assign cosLUT_MPORT_523_en = reset;
  assign cosLUT_MPORT_524_data = 32'h3f319eda;
  assign cosLUT_MPORT_524_addr = 11'h20c;
  assign cosLUT_MPORT_524_mask = 1'h1;
  assign cosLUT_MPORT_524_en = reset;
  assign cosLUT_MPORT_525_data = 32'h3f315662;
  assign cosLUT_MPORT_525_addr = 11'h20d;
  assign cosLUT_MPORT_525_mask = 1'h1;
  assign cosLUT_MPORT_525_en = reset;
  assign cosLUT_MPORT_526_data = 32'h3f310dcf;
  assign cosLUT_MPORT_526_addr = 11'h20e;
  assign cosLUT_MPORT_526_mask = 1'h1;
  assign cosLUT_MPORT_526_en = reset;
  assign cosLUT_MPORT_527_data = 32'h3f30c521;
  assign cosLUT_MPORT_527_addr = 11'h20f;
  assign cosLUT_MPORT_527_mask = 1'h1;
  assign cosLUT_MPORT_527_en = reset;
  assign cosLUT_MPORT_528_data = 32'h3f307c57;
  assign cosLUT_MPORT_528_addr = 11'h210;
  assign cosLUT_MPORT_528_mask = 1'h1;
  assign cosLUT_MPORT_528_en = reset;
  assign cosLUT_MPORT_529_data = 32'h3f303372;
  assign cosLUT_MPORT_529_addr = 11'h211;
  assign cosLUT_MPORT_529_mask = 1'h1;
  assign cosLUT_MPORT_529_en = reset;
  assign cosLUT_MPORT_530_data = 32'h3f2fea72;
  assign cosLUT_MPORT_530_addr = 11'h212;
  assign cosLUT_MPORT_530_mask = 1'h1;
  assign cosLUT_MPORT_530_en = reset;
  assign cosLUT_MPORT_531_data = 32'h3f2fa157;
  assign cosLUT_MPORT_531_addr = 11'h213;
  assign cosLUT_MPORT_531_mask = 1'h1;
  assign cosLUT_MPORT_531_en = reset;
  assign cosLUT_MPORT_532_data = 32'h3f2f5821;
  assign cosLUT_MPORT_532_addr = 11'h214;
  assign cosLUT_MPORT_532_mask = 1'h1;
  assign cosLUT_MPORT_532_en = reset;
  assign cosLUT_MPORT_533_data = 32'h3f2f0ed0;
  assign cosLUT_MPORT_533_addr = 11'h215;
  assign cosLUT_MPORT_533_mask = 1'h1;
  assign cosLUT_MPORT_533_en = reset;
  assign cosLUT_MPORT_534_data = 32'h3f2ec563;
  assign cosLUT_MPORT_534_addr = 11'h216;
  assign cosLUT_MPORT_534_mask = 1'h1;
  assign cosLUT_MPORT_534_en = reset;
  assign cosLUT_MPORT_535_data = 32'h3f2e7bdc;
  assign cosLUT_MPORT_535_addr = 11'h217;
  assign cosLUT_MPORT_535_mask = 1'h1;
  assign cosLUT_MPORT_535_en = reset;
  assign cosLUT_MPORT_536_data = 32'h3f2e323a;
  assign cosLUT_MPORT_536_addr = 11'h218;
  assign cosLUT_MPORT_536_mask = 1'h1;
  assign cosLUT_MPORT_536_en = reset;
  assign cosLUT_MPORT_537_data = 32'h3f2de87d;
  assign cosLUT_MPORT_537_addr = 11'h219;
  assign cosLUT_MPORT_537_mask = 1'h1;
  assign cosLUT_MPORT_537_en = reset;
  assign cosLUT_MPORT_538_data = 32'h3f2d9ea5;
  assign cosLUT_MPORT_538_addr = 11'h21a;
  assign cosLUT_MPORT_538_mask = 1'h1;
  assign cosLUT_MPORT_538_en = reset;
  assign cosLUT_MPORT_539_data = 32'h3f2d54b2;
  assign cosLUT_MPORT_539_addr = 11'h21b;
  assign cosLUT_MPORT_539_mask = 1'h1;
  assign cosLUT_MPORT_539_en = reset;
  assign cosLUT_MPORT_540_data = 32'h3f2d0aa5;
  assign cosLUT_MPORT_540_addr = 11'h21c;
  assign cosLUT_MPORT_540_mask = 1'h1;
  assign cosLUT_MPORT_540_en = reset;
  assign cosLUT_MPORT_541_data = 32'h3f2cc07c;
  assign cosLUT_MPORT_541_addr = 11'h21d;
  assign cosLUT_MPORT_541_mask = 1'h1;
  assign cosLUT_MPORT_541_en = reset;
  assign cosLUT_MPORT_542_data = 32'h3f2c763a;
  assign cosLUT_MPORT_542_addr = 11'h21e;
  assign cosLUT_MPORT_542_mask = 1'h1;
  assign cosLUT_MPORT_542_en = reset;
  assign cosLUT_MPORT_543_data = 32'h3f2c2bdc;
  assign cosLUT_MPORT_543_addr = 11'h21f;
  assign cosLUT_MPORT_543_mask = 1'h1;
  assign cosLUT_MPORT_543_en = reset;
  assign cosLUT_MPORT_544_data = 32'h3f2be164;
  assign cosLUT_MPORT_544_addr = 11'h220;
  assign cosLUT_MPORT_544_mask = 1'h1;
  assign cosLUT_MPORT_544_en = reset;
  assign cosLUT_MPORT_545_data = 32'h3f2b96d2;
  assign cosLUT_MPORT_545_addr = 11'h221;
  assign cosLUT_MPORT_545_mask = 1'h1;
  assign cosLUT_MPORT_545_en = reset;
  assign cosLUT_MPORT_546_data = 32'h3f2b4c25;
  assign cosLUT_MPORT_546_addr = 11'h222;
  assign cosLUT_MPORT_546_mask = 1'h1;
  assign cosLUT_MPORT_546_en = reset;
  assign cosLUT_MPORT_547_data = 32'h3f2b015d;
  assign cosLUT_MPORT_547_addr = 11'h223;
  assign cosLUT_MPORT_547_mask = 1'h1;
  assign cosLUT_MPORT_547_en = reset;
  assign cosLUT_MPORT_548_data = 32'h3f2ab67c;
  assign cosLUT_MPORT_548_addr = 11'h224;
  assign cosLUT_MPORT_548_mask = 1'h1;
  assign cosLUT_MPORT_548_en = reset;
  assign cosLUT_MPORT_549_data = 32'h3f2a6b7f;
  assign cosLUT_MPORT_549_addr = 11'h225;
  assign cosLUT_MPORT_549_mask = 1'h1;
  assign cosLUT_MPORT_549_en = reset;
  assign cosLUT_MPORT_550_data = 32'h3f2a2069;
  assign cosLUT_MPORT_550_addr = 11'h226;
  assign cosLUT_MPORT_550_mask = 1'h1;
  assign cosLUT_MPORT_550_en = reset;
  assign cosLUT_MPORT_551_data = 32'h3f29d538;
  assign cosLUT_MPORT_551_addr = 11'h227;
  assign cosLUT_MPORT_551_mask = 1'h1;
  assign cosLUT_MPORT_551_en = reset;
  assign cosLUT_MPORT_552_data = 32'h3f2989ed;
  assign cosLUT_MPORT_552_addr = 11'h228;
  assign cosLUT_MPORT_552_mask = 1'h1;
  assign cosLUT_MPORT_552_en = reset;
  assign cosLUT_MPORT_553_data = 32'h3f293e88;
  assign cosLUT_MPORT_553_addr = 11'h229;
  assign cosLUT_MPORT_553_mask = 1'h1;
  assign cosLUT_MPORT_553_en = reset;
  assign cosLUT_MPORT_554_data = 32'h3f28f309;
  assign cosLUT_MPORT_554_addr = 11'h22a;
  assign cosLUT_MPORT_554_mask = 1'h1;
  assign cosLUT_MPORT_554_en = reset;
  assign cosLUT_MPORT_555_data = 32'h3f28a770;
  assign cosLUT_MPORT_555_addr = 11'h22b;
  assign cosLUT_MPORT_555_mask = 1'h1;
  assign cosLUT_MPORT_555_en = reset;
  assign cosLUT_MPORT_556_data = 32'h3f285bbd;
  assign cosLUT_MPORT_556_addr = 11'h22c;
  assign cosLUT_MPORT_556_mask = 1'h1;
  assign cosLUT_MPORT_556_en = reset;
  assign cosLUT_MPORT_557_data = 32'h3f280ff0;
  assign cosLUT_MPORT_557_addr = 11'h22d;
  assign cosLUT_MPORT_557_mask = 1'h1;
  assign cosLUT_MPORT_557_en = reset;
  assign cosLUT_MPORT_558_data = 32'h3f27c409;
  assign cosLUT_MPORT_558_addr = 11'h22e;
  assign cosLUT_MPORT_558_mask = 1'h1;
  assign cosLUT_MPORT_558_en = reset;
  assign cosLUT_MPORT_559_data = 32'h3f277808;
  assign cosLUT_MPORT_559_addr = 11'h22f;
  assign cosLUT_MPORT_559_mask = 1'h1;
  assign cosLUT_MPORT_559_en = reset;
  assign cosLUT_MPORT_560_data = 32'h3f272bed;
  assign cosLUT_MPORT_560_addr = 11'h230;
  assign cosLUT_MPORT_560_mask = 1'h1;
  assign cosLUT_MPORT_560_en = reset;
  assign cosLUT_MPORT_561_data = 32'h3f26dfb8;
  assign cosLUT_MPORT_561_addr = 11'h231;
  assign cosLUT_MPORT_561_mask = 1'h1;
  assign cosLUT_MPORT_561_en = reset;
  assign cosLUT_MPORT_562_data = 32'h3f26936a;
  assign cosLUT_MPORT_562_addr = 11'h232;
  assign cosLUT_MPORT_562_mask = 1'h1;
  assign cosLUT_MPORT_562_en = reset;
  assign cosLUT_MPORT_563_data = 32'h3f264702;
  assign cosLUT_MPORT_563_addr = 11'h233;
  assign cosLUT_MPORT_563_mask = 1'h1;
  assign cosLUT_MPORT_563_en = reset;
  assign cosLUT_MPORT_564_data = 32'h3f25fa80;
  assign cosLUT_MPORT_564_addr = 11'h234;
  assign cosLUT_MPORT_564_mask = 1'h1;
  assign cosLUT_MPORT_564_en = reset;
  assign cosLUT_MPORT_565_data = 32'h3f25ade4;
  assign cosLUT_MPORT_565_addr = 11'h235;
  assign cosLUT_MPORT_565_mask = 1'h1;
  assign cosLUT_MPORT_565_en = reset;
  assign cosLUT_MPORT_566_data = 32'h3f256130;
  assign cosLUT_MPORT_566_addr = 11'h236;
  assign cosLUT_MPORT_566_mask = 1'h1;
  assign cosLUT_MPORT_566_en = reset;
  assign cosLUT_MPORT_567_data = 32'h3f251461;
  assign cosLUT_MPORT_567_addr = 11'h237;
  assign cosLUT_MPORT_567_mask = 1'h1;
  assign cosLUT_MPORT_567_en = reset;
  assign cosLUT_MPORT_568_data = 32'h3f24c779;
  assign cosLUT_MPORT_568_addr = 11'h238;
  assign cosLUT_MPORT_568_mask = 1'h1;
  assign cosLUT_MPORT_568_en = reset;
  assign cosLUT_MPORT_569_data = 32'h3f247a78;
  assign cosLUT_MPORT_569_addr = 11'h239;
  assign cosLUT_MPORT_569_mask = 1'h1;
  assign cosLUT_MPORT_569_en = reset;
  assign cosLUT_MPORT_570_data = 32'h3f242d5d;
  assign cosLUT_MPORT_570_addr = 11'h23a;
  assign cosLUT_MPORT_570_mask = 1'h1;
  assign cosLUT_MPORT_570_en = reset;
  assign cosLUT_MPORT_571_data = 32'h3f23e029;
  assign cosLUT_MPORT_571_addr = 11'h23b;
  assign cosLUT_MPORT_571_mask = 1'h1;
  assign cosLUT_MPORT_571_en = reset;
  assign cosLUT_MPORT_572_data = 32'h3f2392dc;
  assign cosLUT_MPORT_572_addr = 11'h23c;
  assign cosLUT_MPORT_572_mask = 1'h1;
  assign cosLUT_MPORT_572_en = reset;
  assign cosLUT_MPORT_573_data = 32'h3f234575;
  assign cosLUT_MPORT_573_addr = 11'h23d;
  assign cosLUT_MPORT_573_mask = 1'h1;
  assign cosLUT_MPORT_573_en = reset;
  assign cosLUT_MPORT_574_data = 32'h3f22f7f5;
  assign cosLUT_MPORT_574_addr = 11'h23e;
  assign cosLUT_MPORT_574_mask = 1'h1;
  assign cosLUT_MPORT_574_en = reset;
  assign cosLUT_MPORT_575_data = 32'h3f22aa5d;
  assign cosLUT_MPORT_575_addr = 11'h23f;
  assign cosLUT_MPORT_575_mask = 1'h1;
  assign cosLUT_MPORT_575_en = reset;
  assign cosLUT_MPORT_576_data = 32'h3f225cab;
  assign cosLUT_MPORT_576_addr = 11'h240;
  assign cosLUT_MPORT_576_mask = 1'h1;
  assign cosLUT_MPORT_576_en = reset;
  assign cosLUT_MPORT_577_data = 32'h3f220ee0;
  assign cosLUT_MPORT_577_addr = 11'h241;
  assign cosLUT_MPORT_577_mask = 1'h1;
  assign cosLUT_MPORT_577_en = reset;
  assign cosLUT_MPORT_578_data = 32'h3f21c0fc;
  assign cosLUT_MPORT_578_addr = 11'h242;
  assign cosLUT_MPORT_578_mask = 1'h1;
  assign cosLUT_MPORT_578_en = reset;
  assign cosLUT_MPORT_579_data = 32'h3f2172ff;
  assign cosLUT_MPORT_579_addr = 11'h243;
  assign cosLUT_MPORT_579_mask = 1'h1;
  assign cosLUT_MPORT_579_en = reset;
  assign cosLUT_MPORT_580_data = 32'h3f2124e9;
  assign cosLUT_MPORT_580_addr = 11'h244;
  assign cosLUT_MPORT_580_mask = 1'h1;
  assign cosLUT_MPORT_580_en = reset;
  assign cosLUT_MPORT_581_data = 32'h3f20d6ba;
  assign cosLUT_MPORT_581_addr = 11'h245;
  assign cosLUT_MPORT_581_mask = 1'h1;
  assign cosLUT_MPORT_581_en = reset;
  assign cosLUT_MPORT_582_data = 32'h3f208872;
  assign cosLUT_MPORT_582_addr = 11'h246;
  assign cosLUT_MPORT_582_mask = 1'h1;
  assign cosLUT_MPORT_582_en = reset;
  assign cosLUT_MPORT_583_data = 32'h3f203a12;
  assign cosLUT_MPORT_583_addr = 11'h247;
  assign cosLUT_MPORT_583_mask = 1'h1;
  assign cosLUT_MPORT_583_en = reset;
  assign cosLUT_MPORT_584_data = 32'h3f1feb99;
  assign cosLUT_MPORT_584_addr = 11'h248;
  assign cosLUT_MPORT_584_mask = 1'h1;
  assign cosLUT_MPORT_584_en = reset;
  assign cosLUT_MPORT_585_data = 32'h3f1f9d07;
  assign cosLUT_MPORT_585_addr = 11'h249;
  assign cosLUT_MPORT_585_mask = 1'h1;
  assign cosLUT_MPORT_585_en = reset;
  assign cosLUT_MPORT_586_data = 32'h3f1f4e5d;
  assign cosLUT_MPORT_586_addr = 11'h24a;
  assign cosLUT_MPORT_586_mask = 1'h1;
  assign cosLUT_MPORT_586_en = reset;
  assign cosLUT_MPORT_587_data = 32'h3f1eff9a;
  assign cosLUT_MPORT_587_addr = 11'h24b;
  assign cosLUT_MPORT_587_mask = 1'h1;
  assign cosLUT_MPORT_587_en = reset;
  assign cosLUT_MPORT_588_data = 32'h3f1eb0be;
  assign cosLUT_MPORT_588_addr = 11'h24c;
  assign cosLUT_MPORT_588_mask = 1'h1;
  assign cosLUT_MPORT_588_en = reset;
  assign cosLUT_MPORT_589_data = 32'h3f1e61ca;
  assign cosLUT_MPORT_589_addr = 11'h24d;
  assign cosLUT_MPORT_589_mask = 1'h1;
  assign cosLUT_MPORT_589_en = reset;
  assign cosLUT_MPORT_590_data = 32'h3f1e12be;
  assign cosLUT_MPORT_590_addr = 11'h24e;
  assign cosLUT_MPORT_590_mask = 1'h1;
  assign cosLUT_MPORT_590_en = reset;
  assign cosLUT_MPORT_591_data = 32'h3f1dc399;
  assign cosLUT_MPORT_591_addr = 11'h24f;
  assign cosLUT_MPORT_591_mask = 1'h1;
  assign cosLUT_MPORT_591_en = reset;
  assign cosLUT_MPORT_592_data = 32'h3f1d745c;
  assign cosLUT_MPORT_592_addr = 11'h250;
  assign cosLUT_MPORT_592_mask = 1'h1;
  assign cosLUT_MPORT_592_en = reset;
  assign cosLUT_MPORT_593_data = 32'h3f1d2507;
  assign cosLUT_MPORT_593_addr = 11'h251;
  assign cosLUT_MPORT_593_mask = 1'h1;
  assign cosLUT_MPORT_593_en = reset;
  assign cosLUT_MPORT_594_data = 32'h3f1cd599;
  assign cosLUT_MPORT_594_addr = 11'h252;
  assign cosLUT_MPORT_594_mask = 1'h1;
  assign cosLUT_MPORT_594_en = reset;
  assign cosLUT_MPORT_595_data = 32'h3f1c8613;
  assign cosLUT_MPORT_595_addr = 11'h253;
  assign cosLUT_MPORT_595_mask = 1'h1;
  assign cosLUT_MPORT_595_en = reset;
  assign cosLUT_MPORT_596_data = 32'h3f1c3675;
  assign cosLUT_MPORT_596_addr = 11'h254;
  assign cosLUT_MPORT_596_mask = 1'h1;
  assign cosLUT_MPORT_596_en = reset;
  assign cosLUT_MPORT_597_data = 32'h3f1be6bf;
  assign cosLUT_MPORT_597_addr = 11'h255;
  assign cosLUT_MPORT_597_mask = 1'h1;
  assign cosLUT_MPORT_597_en = reset;
  assign cosLUT_MPORT_598_data = 32'h3f1b96f1;
  assign cosLUT_MPORT_598_addr = 11'h256;
  assign cosLUT_MPORT_598_mask = 1'h1;
  assign cosLUT_MPORT_598_en = reset;
  assign cosLUT_MPORT_599_data = 32'h3f1b470a;
  assign cosLUT_MPORT_599_addr = 11'h257;
  assign cosLUT_MPORT_599_mask = 1'h1;
  assign cosLUT_MPORT_599_en = reset;
  assign cosLUT_MPORT_600_data = 32'h3f1af70c;
  assign cosLUT_MPORT_600_addr = 11'h258;
  assign cosLUT_MPORT_600_mask = 1'h1;
  assign cosLUT_MPORT_600_en = reset;
  assign cosLUT_MPORT_601_data = 32'h3f1aa6f6;
  assign cosLUT_MPORT_601_addr = 11'h259;
  assign cosLUT_MPORT_601_mask = 1'h1;
  assign cosLUT_MPORT_601_en = reset;
  assign cosLUT_MPORT_602_data = 32'h3f1a56c8;
  assign cosLUT_MPORT_602_addr = 11'h25a;
  assign cosLUT_MPORT_602_mask = 1'h1;
  assign cosLUT_MPORT_602_en = reset;
  assign cosLUT_MPORT_603_data = 32'h3f1a0683;
  assign cosLUT_MPORT_603_addr = 11'h25b;
  assign cosLUT_MPORT_603_mask = 1'h1;
  assign cosLUT_MPORT_603_en = reset;
  assign cosLUT_MPORT_604_data = 32'h3f19b625;
  assign cosLUT_MPORT_604_addr = 11'h25c;
  assign cosLUT_MPORT_604_mask = 1'h1;
  assign cosLUT_MPORT_604_en = reset;
  assign cosLUT_MPORT_605_data = 32'h3f1965b0;
  assign cosLUT_MPORT_605_addr = 11'h25d;
  assign cosLUT_MPORT_605_mask = 1'h1;
  assign cosLUT_MPORT_605_en = reset;
  assign cosLUT_MPORT_606_data = 32'h3f191523;
  assign cosLUT_MPORT_606_addr = 11'h25e;
  assign cosLUT_MPORT_606_mask = 1'h1;
  assign cosLUT_MPORT_606_en = reset;
  assign cosLUT_MPORT_607_data = 32'h3f18c47f;
  assign cosLUT_MPORT_607_addr = 11'h25f;
  assign cosLUT_MPORT_607_mask = 1'h1;
  assign cosLUT_MPORT_607_en = reset;
  assign cosLUT_MPORT_608_data = 32'h3f1873c2;
  assign cosLUT_MPORT_608_addr = 11'h260;
  assign cosLUT_MPORT_608_mask = 1'h1;
  assign cosLUT_MPORT_608_en = reset;
  assign cosLUT_MPORT_609_data = 32'h3f1822ef;
  assign cosLUT_MPORT_609_addr = 11'h261;
  assign cosLUT_MPORT_609_mask = 1'h1;
  assign cosLUT_MPORT_609_en = reset;
  assign cosLUT_MPORT_610_data = 32'h3f17d204;
  assign cosLUT_MPORT_610_addr = 11'h262;
  assign cosLUT_MPORT_610_mask = 1'h1;
  assign cosLUT_MPORT_610_en = reset;
  assign cosLUT_MPORT_611_data = 32'h3f178101;
  assign cosLUT_MPORT_611_addr = 11'h263;
  assign cosLUT_MPORT_611_mask = 1'h1;
  assign cosLUT_MPORT_611_en = reset;
  assign cosLUT_MPORT_612_data = 32'h3f172fe8;
  assign cosLUT_MPORT_612_addr = 11'h264;
  assign cosLUT_MPORT_612_mask = 1'h1;
  assign cosLUT_MPORT_612_en = reset;
  assign cosLUT_MPORT_613_data = 32'h3f16deb6;
  assign cosLUT_MPORT_613_addr = 11'h265;
  assign cosLUT_MPORT_613_mask = 1'h1;
  assign cosLUT_MPORT_613_en = reset;
  assign cosLUT_MPORT_614_data = 32'h3f168d6e;
  assign cosLUT_MPORT_614_addr = 11'h266;
  assign cosLUT_MPORT_614_mask = 1'h1;
  assign cosLUT_MPORT_614_en = reset;
  assign cosLUT_MPORT_615_data = 32'h3f163c0e;
  assign cosLUT_MPORT_615_addr = 11'h267;
  assign cosLUT_MPORT_615_mask = 1'h1;
  assign cosLUT_MPORT_615_en = reset;
  assign cosLUT_MPORT_616_data = 32'h3f15ea97;
  assign cosLUT_MPORT_616_addr = 11'h268;
  assign cosLUT_MPORT_616_mask = 1'h1;
  assign cosLUT_MPORT_616_en = reset;
  assign cosLUT_MPORT_617_data = 32'h3f159909;
  assign cosLUT_MPORT_617_addr = 11'h269;
  assign cosLUT_MPORT_617_mask = 1'h1;
  assign cosLUT_MPORT_617_en = reset;
  assign cosLUT_MPORT_618_data = 32'h3f154764;
  assign cosLUT_MPORT_618_addr = 11'h26a;
  assign cosLUT_MPORT_618_mask = 1'h1;
  assign cosLUT_MPORT_618_en = reset;
  assign cosLUT_MPORT_619_data = 32'h3f14f5a8;
  assign cosLUT_MPORT_619_addr = 11'h26b;
  assign cosLUT_MPORT_619_mask = 1'h1;
  assign cosLUT_MPORT_619_en = reset;
  assign cosLUT_MPORT_620_data = 32'h3f14a3d5;
  assign cosLUT_MPORT_620_addr = 11'h26c;
  assign cosLUT_MPORT_620_mask = 1'h1;
  assign cosLUT_MPORT_620_en = reset;
  assign cosLUT_MPORT_621_data = 32'h3f1451eb;
  assign cosLUT_MPORT_621_addr = 11'h26d;
  assign cosLUT_MPORT_621_mask = 1'h1;
  assign cosLUT_MPORT_621_en = reset;
  assign cosLUT_MPORT_622_data = 32'h3f13ffea;
  assign cosLUT_MPORT_622_addr = 11'h26e;
  assign cosLUT_MPORT_622_mask = 1'h1;
  assign cosLUT_MPORT_622_en = reset;
  assign cosLUT_MPORT_623_data = 32'h3f13add2;
  assign cosLUT_MPORT_623_addr = 11'h26f;
  assign cosLUT_MPORT_623_mask = 1'h1;
  assign cosLUT_MPORT_623_en = reset;
  assign cosLUT_MPORT_624_data = 32'h3f135ba4;
  assign cosLUT_MPORT_624_addr = 11'h270;
  assign cosLUT_MPORT_624_mask = 1'h1;
  assign cosLUT_MPORT_624_en = reset;
  assign cosLUT_MPORT_625_data = 32'h3f13095f;
  assign cosLUT_MPORT_625_addr = 11'h271;
  assign cosLUT_MPORT_625_mask = 1'h1;
  assign cosLUT_MPORT_625_en = reset;
  assign cosLUT_MPORT_626_data = 32'h3f12b703;
  assign cosLUT_MPORT_626_addr = 11'h272;
  assign cosLUT_MPORT_626_mask = 1'h1;
  assign cosLUT_MPORT_626_en = reset;
  assign cosLUT_MPORT_627_data = 32'h3f126490;
  assign cosLUT_MPORT_627_addr = 11'h273;
  assign cosLUT_MPORT_627_mask = 1'h1;
  assign cosLUT_MPORT_627_en = reset;
  assign cosLUT_MPORT_628_data = 32'h3f121207;
  assign cosLUT_MPORT_628_addr = 11'h274;
  assign cosLUT_MPORT_628_mask = 1'h1;
  assign cosLUT_MPORT_628_en = reset;
  assign cosLUT_MPORT_629_data = 32'h3f11bf67;
  assign cosLUT_MPORT_629_addr = 11'h275;
  assign cosLUT_MPORT_629_mask = 1'h1;
  assign cosLUT_MPORT_629_en = reset;
  assign cosLUT_MPORT_630_data = 32'h3f116cb1;
  assign cosLUT_MPORT_630_addr = 11'h276;
  assign cosLUT_MPORT_630_mask = 1'h1;
  assign cosLUT_MPORT_630_en = reset;
  assign cosLUT_MPORT_631_data = 32'h3f1119e4;
  assign cosLUT_MPORT_631_addr = 11'h277;
  assign cosLUT_MPORT_631_mask = 1'h1;
  assign cosLUT_MPORT_631_en = reset;
  assign cosLUT_MPORT_632_data = 32'h3f10c701;
  assign cosLUT_MPORT_632_addr = 11'h278;
  assign cosLUT_MPORT_632_mask = 1'h1;
  assign cosLUT_MPORT_632_en = reset;
  assign cosLUT_MPORT_633_data = 32'h3f107408;
  assign cosLUT_MPORT_633_addr = 11'h279;
  assign cosLUT_MPORT_633_mask = 1'h1;
  assign cosLUT_MPORT_633_en = reset;
  assign cosLUT_MPORT_634_data = 32'h3f1020f8;
  assign cosLUT_MPORT_634_addr = 11'h27a;
  assign cosLUT_MPORT_634_mask = 1'h1;
  assign cosLUT_MPORT_634_en = reset;
  assign cosLUT_MPORT_635_data = 32'h3f0fcdd2;
  assign cosLUT_MPORT_635_addr = 11'h27b;
  assign cosLUT_MPORT_635_mask = 1'h1;
  assign cosLUT_MPORT_635_en = reset;
  assign cosLUT_MPORT_636_data = 32'h3f0f7a96;
  assign cosLUT_MPORT_636_addr = 11'h27c;
  assign cosLUT_MPORT_636_mask = 1'h1;
  assign cosLUT_MPORT_636_en = reset;
  assign cosLUT_MPORT_637_data = 32'h3f0f2744;
  assign cosLUT_MPORT_637_addr = 11'h27d;
  assign cosLUT_MPORT_637_mask = 1'h1;
  assign cosLUT_MPORT_637_en = reset;
  assign cosLUT_MPORT_638_data = 32'h3f0ed3dc;
  assign cosLUT_MPORT_638_addr = 11'h27e;
  assign cosLUT_MPORT_638_mask = 1'h1;
  assign cosLUT_MPORT_638_en = reset;
  assign cosLUT_MPORT_639_data = 32'h3f0e805d;
  assign cosLUT_MPORT_639_addr = 11'h27f;
  assign cosLUT_MPORT_639_mask = 1'h1;
  assign cosLUT_MPORT_639_en = reset;
  assign cosLUT_MPORT_640_data = 32'h3f0e2cc9;
  assign cosLUT_MPORT_640_addr = 11'h280;
  assign cosLUT_MPORT_640_mask = 1'h1;
  assign cosLUT_MPORT_640_en = reset;
  assign cosLUT_MPORT_641_data = 32'h3f0dd91f;
  assign cosLUT_MPORT_641_addr = 11'h281;
  assign cosLUT_MPORT_641_mask = 1'h1;
  assign cosLUT_MPORT_641_en = reset;
  assign cosLUT_MPORT_642_data = 32'h3f0d855f;
  assign cosLUT_MPORT_642_addr = 11'h282;
  assign cosLUT_MPORT_642_mask = 1'h1;
  assign cosLUT_MPORT_642_en = reset;
  assign cosLUT_MPORT_643_data = 32'h3f0d3189;
  assign cosLUT_MPORT_643_addr = 11'h283;
  assign cosLUT_MPORT_643_mask = 1'h1;
  assign cosLUT_MPORT_643_en = reset;
  assign cosLUT_MPORT_644_data = 32'h3f0cdd9d;
  assign cosLUT_MPORT_644_addr = 11'h284;
  assign cosLUT_MPORT_644_mask = 1'h1;
  assign cosLUT_MPORT_644_en = reset;
  assign cosLUT_MPORT_645_data = 32'h3f0c899c;
  assign cosLUT_MPORT_645_addr = 11'h285;
  assign cosLUT_MPORT_645_mask = 1'h1;
  assign cosLUT_MPORT_645_en = reset;
  assign cosLUT_MPORT_646_data = 32'h3f0c3584;
  assign cosLUT_MPORT_646_addr = 11'h286;
  assign cosLUT_MPORT_646_mask = 1'h1;
  assign cosLUT_MPORT_646_en = reset;
  assign cosLUT_MPORT_647_data = 32'h3f0be158;
  assign cosLUT_MPORT_647_addr = 11'h287;
  assign cosLUT_MPORT_647_mask = 1'h1;
  assign cosLUT_MPORT_647_en = reset;
  assign cosLUT_MPORT_648_data = 32'h3f0b8d15;
  assign cosLUT_MPORT_648_addr = 11'h288;
  assign cosLUT_MPORT_648_mask = 1'h1;
  assign cosLUT_MPORT_648_en = reset;
  assign cosLUT_MPORT_649_data = 32'h3f0b38bd;
  assign cosLUT_MPORT_649_addr = 11'h289;
  assign cosLUT_MPORT_649_mask = 1'h1;
  assign cosLUT_MPORT_649_en = reset;
  assign cosLUT_MPORT_650_data = 32'h3f0ae450;
  assign cosLUT_MPORT_650_addr = 11'h28a;
  assign cosLUT_MPORT_650_mask = 1'h1;
  assign cosLUT_MPORT_650_en = reset;
  assign cosLUT_MPORT_651_data = 32'h3f0a8fcd;
  assign cosLUT_MPORT_651_addr = 11'h28b;
  assign cosLUT_MPORT_651_mask = 1'h1;
  assign cosLUT_MPORT_651_en = reset;
  assign cosLUT_MPORT_652_data = 32'h3f0a3b35;
  assign cosLUT_MPORT_652_addr = 11'h28c;
  assign cosLUT_MPORT_652_mask = 1'h1;
  assign cosLUT_MPORT_652_en = reset;
  assign cosLUT_MPORT_653_data = 32'h3f09e687;
  assign cosLUT_MPORT_653_addr = 11'h28d;
  assign cosLUT_MPORT_653_mask = 1'h1;
  assign cosLUT_MPORT_653_en = reset;
  assign cosLUT_MPORT_654_data = 32'h3f0991c4;
  assign cosLUT_MPORT_654_addr = 11'h28e;
  assign cosLUT_MPORT_654_mask = 1'h1;
  assign cosLUT_MPORT_654_en = reset;
  assign cosLUT_MPORT_655_data = 32'h3f093cec;
  assign cosLUT_MPORT_655_addr = 11'h28f;
  assign cosLUT_MPORT_655_mask = 1'h1;
  assign cosLUT_MPORT_655_en = reset;
  assign cosLUT_MPORT_656_data = 32'h3f08e7ff;
  assign cosLUT_MPORT_656_addr = 11'h290;
  assign cosLUT_MPORT_656_mask = 1'h1;
  assign cosLUT_MPORT_656_en = reset;
  assign cosLUT_MPORT_657_data = 32'h3f0892fd;
  assign cosLUT_MPORT_657_addr = 11'h291;
  assign cosLUT_MPORT_657_mask = 1'h1;
  assign cosLUT_MPORT_657_en = reset;
  assign cosLUT_MPORT_658_data = 32'h3f083de5;
  assign cosLUT_MPORT_658_addr = 11'h292;
  assign cosLUT_MPORT_658_mask = 1'h1;
  assign cosLUT_MPORT_658_en = reset;
  assign cosLUT_MPORT_659_data = 32'h3f07e8b9;
  assign cosLUT_MPORT_659_addr = 11'h293;
  assign cosLUT_MPORT_659_mask = 1'h1;
  assign cosLUT_MPORT_659_en = reset;
  assign cosLUT_MPORT_660_data = 32'h3f079378;
  assign cosLUT_MPORT_660_addr = 11'h294;
  assign cosLUT_MPORT_660_mask = 1'h1;
  assign cosLUT_MPORT_660_en = reset;
  assign cosLUT_MPORT_661_data = 32'h3f073e21;
  assign cosLUT_MPORT_661_addr = 11'h295;
  assign cosLUT_MPORT_661_mask = 1'h1;
  assign cosLUT_MPORT_661_en = reset;
  assign cosLUT_MPORT_662_data = 32'h3f06e8b6;
  assign cosLUT_MPORT_662_addr = 11'h296;
  assign cosLUT_MPORT_662_mask = 1'h1;
  assign cosLUT_MPORT_662_en = reset;
  assign cosLUT_MPORT_663_data = 32'h3f069336;
  assign cosLUT_MPORT_663_addr = 11'h297;
  assign cosLUT_MPORT_663_mask = 1'h1;
  assign cosLUT_MPORT_663_en = reset;
  assign cosLUT_MPORT_664_data = 32'h3f063da1;
  assign cosLUT_MPORT_664_addr = 11'h298;
  assign cosLUT_MPORT_664_mask = 1'h1;
  assign cosLUT_MPORT_664_en = reset;
  assign cosLUT_MPORT_665_data = 32'h3f05e7f8;
  assign cosLUT_MPORT_665_addr = 11'h299;
  assign cosLUT_MPORT_665_mask = 1'h1;
  assign cosLUT_MPORT_665_en = reset;
  assign cosLUT_MPORT_666_data = 32'h3f05923a;
  assign cosLUT_MPORT_666_addr = 11'h29a;
  assign cosLUT_MPORT_666_mask = 1'h1;
  assign cosLUT_MPORT_666_en = reset;
  assign cosLUT_MPORT_667_data = 32'h3f053c67;
  assign cosLUT_MPORT_667_addr = 11'h29b;
  assign cosLUT_MPORT_667_mask = 1'h1;
  assign cosLUT_MPORT_667_en = reset;
  assign cosLUT_MPORT_668_data = 32'h3f04e680;
  assign cosLUT_MPORT_668_addr = 11'h29c;
  assign cosLUT_MPORT_668_mask = 1'h1;
  assign cosLUT_MPORT_668_en = reset;
  assign cosLUT_MPORT_669_data = 32'h3f049084;
  assign cosLUT_MPORT_669_addr = 11'h29d;
  assign cosLUT_MPORT_669_mask = 1'h1;
  assign cosLUT_MPORT_669_en = reset;
  assign cosLUT_MPORT_670_data = 32'h3f043a74;
  assign cosLUT_MPORT_670_addr = 11'h29e;
  assign cosLUT_MPORT_670_mask = 1'h1;
  assign cosLUT_MPORT_670_en = reset;
  assign cosLUT_MPORT_671_data = 32'h3f03e44f;
  assign cosLUT_MPORT_671_addr = 11'h29f;
  assign cosLUT_MPORT_671_mask = 1'h1;
  assign cosLUT_MPORT_671_en = reset;
  assign cosLUT_MPORT_672_data = 32'h3f038e16;
  assign cosLUT_MPORT_672_addr = 11'h2a0;
  assign cosLUT_MPORT_672_mask = 1'h1;
  assign cosLUT_MPORT_672_en = reset;
  assign cosLUT_MPORT_673_data = 32'h3f0337c9;
  assign cosLUT_MPORT_673_addr = 11'h2a1;
  assign cosLUT_MPORT_673_mask = 1'h1;
  assign cosLUT_MPORT_673_en = reset;
  assign cosLUT_MPORT_674_data = 32'h3f02e167;
  assign cosLUT_MPORT_674_addr = 11'h2a2;
  assign cosLUT_MPORT_674_mask = 1'h1;
  assign cosLUT_MPORT_674_en = reset;
  assign cosLUT_MPORT_675_data = 32'h3f028af1;
  assign cosLUT_MPORT_675_addr = 11'h2a3;
  assign cosLUT_MPORT_675_mask = 1'h1;
  assign cosLUT_MPORT_675_en = reset;
  assign cosLUT_MPORT_676_data = 32'h3f023468;
  assign cosLUT_MPORT_676_addr = 11'h2a4;
  assign cosLUT_MPORT_676_mask = 1'h1;
  assign cosLUT_MPORT_676_en = reset;
  assign cosLUT_MPORT_677_data = 32'h3f01ddca;
  assign cosLUT_MPORT_677_addr = 11'h2a5;
  assign cosLUT_MPORT_677_mask = 1'h1;
  assign cosLUT_MPORT_677_en = reset;
  assign cosLUT_MPORT_678_data = 32'h3f018718;
  assign cosLUT_MPORT_678_addr = 11'h2a6;
  assign cosLUT_MPORT_678_mask = 1'h1;
  assign cosLUT_MPORT_678_en = reset;
  assign cosLUT_MPORT_679_data = 32'h3f013052;
  assign cosLUT_MPORT_679_addr = 11'h2a7;
  assign cosLUT_MPORT_679_mask = 1'h1;
  assign cosLUT_MPORT_679_en = reset;
  assign cosLUT_MPORT_680_data = 32'h3f00d978;
  assign cosLUT_MPORT_680_addr = 11'h2a8;
  assign cosLUT_MPORT_680_mask = 1'h1;
  assign cosLUT_MPORT_680_en = reset;
  assign cosLUT_MPORT_681_data = 32'h3f00828a;
  assign cosLUT_MPORT_681_addr = 11'h2a9;
  assign cosLUT_MPORT_681_mask = 1'h1;
  assign cosLUT_MPORT_681_en = reset;
  assign cosLUT_MPORT_682_data = 32'h3f002b88;
  assign cosLUT_MPORT_682_addr = 11'h2aa;
  assign cosLUT_MPORT_682_mask = 1'h1;
  assign cosLUT_MPORT_682_en = reset;
  assign cosLUT_MPORT_683_data = 32'h3effa8e6;
  assign cosLUT_MPORT_683_addr = 11'h2ab;
  assign cosLUT_MPORT_683_mask = 1'h1;
  assign cosLUT_MPORT_683_en = reset;
  assign cosLUT_MPORT_684_data = 32'h3efefa93;
  assign cosLUT_MPORT_684_addr = 11'h2ac;
  assign cosLUT_MPORT_684_mask = 1'h1;
  assign cosLUT_MPORT_684_en = reset;
  assign cosLUT_MPORT_685_data = 32'h3efe4c1a;
  assign cosLUT_MPORT_685_addr = 11'h2ad;
  assign cosLUT_MPORT_685_mask = 1'h1;
  assign cosLUT_MPORT_685_en = reset;
  assign cosLUT_MPORT_686_data = 32'h3efd9d79;
  assign cosLUT_MPORT_686_addr = 11'h2ae;
  assign cosLUT_MPORT_686_mask = 1'h1;
  assign cosLUT_MPORT_686_en = reset;
  assign cosLUT_MPORT_687_data = 32'h3efceeb1;
  assign cosLUT_MPORT_687_addr = 11'h2af;
  assign cosLUT_MPORT_687_mask = 1'h1;
  assign cosLUT_MPORT_687_en = reset;
  assign cosLUT_MPORT_688_data = 32'h3efc3fc2;
  assign cosLUT_MPORT_688_addr = 11'h2b0;
  assign cosLUT_MPORT_688_mask = 1'h1;
  assign cosLUT_MPORT_688_en = reset;
  assign cosLUT_MPORT_689_data = 32'h3efb90ac;
  assign cosLUT_MPORT_689_addr = 11'h2b1;
  assign cosLUT_MPORT_689_mask = 1'h1;
  assign cosLUT_MPORT_689_en = reset;
  assign cosLUT_MPORT_690_data = 32'h3efae16f;
  assign cosLUT_MPORT_690_addr = 11'h2b2;
  assign cosLUT_MPORT_690_mask = 1'h1;
  assign cosLUT_MPORT_690_en = reset;
  assign cosLUT_MPORT_691_data = 32'h3efa320c;
  assign cosLUT_MPORT_691_addr = 11'h2b3;
  assign cosLUT_MPORT_691_mask = 1'h1;
  assign cosLUT_MPORT_691_en = reset;
  assign cosLUT_MPORT_692_data = 32'h3ef98282;
  assign cosLUT_MPORT_692_addr = 11'h2b4;
  assign cosLUT_MPORT_692_mask = 1'h1;
  assign cosLUT_MPORT_692_en = reset;
  assign cosLUT_MPORT_693_data = 32'h3ef8d2d1;
  assign cosLUT_MPORT_693_addr = 11'h2b5;
  assign cosLUT_MPORT_693_mask = 1'h1;
  assign cosLUT_MPORT_693_en = reset;
  assign cosLUT_MPORT_694_data = 32'h3ef822fa;
  assign cosLUT_MPORT_694_addr = 11'h2b6;
  assign cosLUT_MPORT_694_mask = 1'h1;
  assign cosLUT_MPORT_694_en = reset;
  assign cosLUT_MPORT_695_data = 32'h3ef772fd;
  assign cosLUT_MPORT_695_addr = 11'h2b7;
  assign cosLUT_MPORT_695_mask = 1'h1;
  assign cosLUT_MPORT_695_en = reset;
  assign cosLUT_MPORT_696_data = 32'h3ef6c2da;
  assign cosLUT_MPORT_696_addr = 11'h2b8;
  assign cosLUT_MPORT_696_mask = 1'h1;
  assign cosLUT_MPORT_696_en = reset;
  assign cosLUT_MPORT_697_data = 32'h3ef61290;
  assign cosLUT_MPORT_697_addr = 11'h2b9;
  assign cosLUT_MPORT_697_mask = 1'h1;
  assign cosLUT_MPORT_697_en = reset;
  assign cosLUT_MPORT_698_data = 32'h3ef56221;
  assign cosLUT_MPORT_698_addr = 11'h2ba;
  assign cosLUT_MPORT_698_mask = 1'h1;
  assign cosLUT_MPORT_698_en = reset;
  assign cosLUT_MPORT_699_data = 32'h3ef4b18c;
  assign cosLUT_MPORT_699_addr = 11'h2bb;
  assign cosLUT_MPORT_699_mask = 1'h1;
  assign cosLUT_MPORT_699_en = reset;
  assign cosLUT_MPORT_700_data = 32'h3ef400d1;
  assign cosLUT_MPORT_700_addr = 11'h2bc;
  assign cosLUT_MPORT_700_mask = 1'h1;
  assign cosLUT_MPORT_700_en = reset;
  assign cosLUT_MPORT_701_data = 32'h3ef34ff0;
  assign cosLUT_MPORT_701_addr = 11'h2bd;
  assign cosLUT_MPORT_701_mask = 1'h1;
  assign cosLUT_MPORT_701_en = reset;
  assign cosLUT_MPORT_702_data = 32'h3ef29eea;
  assign cosLUT_MPORT_702_addr = 11'h2be;
  assign cosLUT_MPORT_702_mask = 1'h1;
  assign cosLUT_MPORT_702_en = reset;
  assign cosLUT_MPORT_703_data = 32'h3ef1edbe;
  assign cosLUT_MPORT_703_addr = 11'h2bf;
  assign cosLUT_MPORT_703_mask = 1'h1;
  assign cosLUT_MPORT_703_en = reset;
  assign cosLUT_MPORT_704_data = 32'h3ef13c6d;
  assign cosLUT_MPORT_704_addr = 11'h2c0;
  assign cosLUT_MPORT_704_mask = 1'h1;
  assign cosLUT_MPORT_704_en = reset;
  assign cosLUT_MPORT_705_data = 32'h3ef08af7;
  assign cosLUT_MPORT_705_addr = 11'h2c1;
  assign cosLUT_MPORT_705_mask = 1'h1;
  assign cosLUT_MPORT_705_en = reset;
  assign cosLUT_MPORT_706_data = 32'h3eefd95c;
  assign cosLUT_MPORT_706_addr = 11'h2c2;
  assign cosLUT_MPORT_706_mask = 1'h1;
  assign cosLUT_MPORT_706_en = reset;
  assign cosLUT_MPORT_707_data = 32'h3eef279b;
  assign cosLUT_MPORT_707_addr = 11'h2c3;
  assign cosLUT_MPORT_707_mask = 1'h1;
  assign cosLUT_MPORT_707_en = reset;
  assign cosLUT_MPORT_708_data = 32'h3eee75b6;
  assign cosLUT_MPORT_708_addr = 11'h2c4;
  assign cosLUT_MPORT_708_mask = 1'h1;
  assign cosLUT_MPORT_708_en = reset;
  assign cosLUT_MPORT_709_data = 32'h3eedc3ac;
  assign cosLUT_MPORT_709_addr = 11'h2c5;
  assign cosLUT_MPORT_709_mask = 1'h1;
  assign cosLUT_MPORT_709_en = reset;
  assign cosLUT_MPORT_710_data = 32'h3eed117d;
  assign cosLUT_MPORT_710_addr = 11'h2c6;
  assign cosLUT_MPORT_710_mask = 1'h1;
  assign cosLUT_MPORT_710_en = reset;
  assign cosLUT_MPORT_711_data = 32'h3eec5f2a;
  assign cosLUT_MPORT_711_addr = 11'h2c7;
  assign cosLUT_MPORT_711_mask = 1'h1;
  assign cosLUT_MPORT_711_en = reset;
  assign cosLUT_MPORT_712_data = 32'h3eebacb2;
  assign cosLUT_MPORT_712_addr = 11'h2c8;
  assign cosLUT_MPORT_712_mask = 1'h1;
  assign cosLUT_MPORT_712_en = reset;
  assign cosLUT_MPORT_713_data = 32'h3eeafa16;
  assign cosLUT_MPORT_713_addr = 11'h2c9;
  assign cosLUT_MPORT_713_mask = 1'h1;
  assign cosLUT_MPORT_713_en = reset;
  assign cosLUT_MPORT_714_data = 32'h3eea4756;
  assign cosLUT_MPORT_714_addr = 11'h2ca;
  assign cosLUT_MPORT_714_mask = 1'h1;
  assign cosLUT_MPORT_714_en = reset;
  assign cosLUT_MPORT_715_data = 32'h3ee99471;
  assign cosLUT_MPORT_715_addr = 11'h2cb;
  assign cosLUT_MPORT_715_mask = 1'h1;
  assign cosLUT_MPORT_715_en = reset;
  assign cosLUT_MPORT_716_data = 32'h3ee8e169;
  assign cosLUT_MPORT_716_addr = 11'h2cc;
  assign cosLUT_MPORT_716_mask = 1'h1;
  assign cosLUT_MPORT_716_en = reset;
  assign cosLUT_MPORT_717_data = 32'h3ee82e3c;
  assign cosLUT_MPORT_717_addr = 11'h2cd;
  assign cosLUT_MPORT_717_mask = 1'h1;
  assign cosLUT_MPORT_717_en = reset;
  assign cosLUT_MPORT_718_data = 32'h3ee77aec;
  assign cosLUT_MPORT_718_addr = 11'h2ce;
  assign cosLUT_MPORT_718_mask = 1'h1;
  assign cosLUT_MPORT_718_en = reset;
  assign cosLUT_MPORT_719_data = 32'h3ee6c778;
  assign cosLUT_MPORT_719_addr = 11'h2cf;
  assign cosLUT_MPORT_719_mask = 1'h1;
  assign cosLUT_MPORT_719_en = reset;
  assign cosLUT_MPORT_720_data = 32'h3ee613e1;
  assign cosLUT_MPORT_720_addr = 11'h2d0;
  assign cosLUT_MPORT_720_mask = 1'h1;
  assign cosLUT_MPORT_720_en = reset;
  assign cosLUT_MPORT_721_data = 32'h3ee56025;
  assign cosLUT_MPORT_721_addr = 11'h2d1;
  assign cosLUT_MPORT_721_mask = 1'h1;
  assign cosLUT_MPORT_721_en = reset;
  assign cosLUT_MPORT_722_data = 32'h3ee4ac47;
  assign cosLUT_MPORT_722_addr = 11'h2d2;
  assign cosLUT_MPORT_722_mask = 1'h1;
  assign cosLUT_MPORT_722_en = reset;
  assign cosLUT_MPORT_723_data = 32'h3ee3f845;
  assign cosLUT_MPORT_723_addr = 11'h2d3;
  assign cosLUT_MPORT_723_mask = 1'h1;
  assign cosLUT_MPORT_723_en = reset;
  assign cosLUT_MPORT_724_data = 32'h3ee34420;
  assign cosLUT_MPORT_724_addr = 11'h2d4;
  assign cosLUT_MPORT_724_mask = 1'h1;
  assign cosLUT_MPORT_724_en = reset;
  assign cosLUT_MPORT_725_data = 32'h3ee28fd8;
  assign cosLUT_MPORT_725_addr = 11'h2d5;
  assign cosLUT_MPORT_725_mask = 1'h1;
  assign cosLUT_MPORT_725_en = reset;
  assign cosLUT_MPORT_726_data = 32'h3ee1db6d;
  assign cosLUT_MPORT_726_addr = 11'h2d6;
  assign cosLUT_MPORT_726_mask = 1'h1;
  assign cosLUT_MPORT_726_en = reset;
  assign cosLUT_MPORT_727_data = 32'h3ee126df;
  assign cosLUT_MPORT_727_addr = 11'h2d7;
  assign cosLUT_MPORT_727_mask = 1'h1;
  assign cosLUT_MPORT_727_en = reset;
  assign cosLUT_MPORT_728_data = 32'h3ee0722f;
  assign cosLUT_MPORT_728_addr = 11'h2d8;
  assign cosLUT_MPORT_728_mask = 1'h1;
  assign cosLUT_MPORT_728_en = reset;
  assign cosLUT_MPORT_729_data = 32'h3edfbd5c;
  assign cosLUT_MPORT_729_addr = 11'h2d9;
  assign cosLUT_MPORT_729_mask = 1'h1;
  assign cosLUT_MPORT_729_en = reset;
  assign cosLUT_MPORT_730_data = 32'h3edf0866;
  assign cosLUT_MPORT_730_addr = 11'h2da;
  assign cosLUT_MPORT_730_mask = 1'h1;
  assign cosLUT_MPORT_730_en = reset;
  assign cosLUT_MPORT_731_data = 32'h3ede534e;
  assign cosLUT_MPORT_731_addr = 11'h2db;
  assign cosLUT_MPORT_731_mask = 1'h1;
  assign cosLUT_MPORT_731_en = reset;
  assign cosLUT_MPORT_732_data = 32'h3edd9e13;
  assign cosLUT_MPORT_732_addr = 11'h2dc;
  assign cosLUT_MPORT_732_mask = 1'h1;
  assign cosLUT_MPORT_732_en = reset;
  assign cosLUT_MPORT_733_data = 32'h3edce8b7;
  assign cosLUT_MPORT_733_addr = 11'h2dd;
  assign cosLUT_MPORT_733_mask = 1'h1;
  assign cosLUT_MPORT_733_en = reset;
  assign cosLUT_MPORT_734_data = 32'h3edc3338;
  assign cosLUT_MPORT_734_addr = 11'h2de;
  assign cosLUT_MPORT_734_mask = 1'h1;
  assign cosLUT_MPORT_734_en = reset;
  assign cosLUT_MPORT_735_data = 32'h3edb7d97;
  assign cosLUT_MPORT_735_addr = 11'h2df;
  assign cosLUT_MPORT_735_mask = 1'h1;
  assign cosLUT_MPORT_735_en = reset;
  assign cosLUT_MPORT_736_data = 32'h3edac7d5;
  assign cosLUT_MPORT_736_addr = 11'h2e0;
  assign cosLUT_MPORT_736_mask = 1'h1;
  assign cosLUT_MPORT_736_en = reset;
  assign cosLUT_MPORT_737_data = 32'h3eda11f1;
  assign cosLUT_MPORT_737_addr = 11'h2e1;
  assign cosLUT_MPORT_737_mask = 1'h1;
  assign cosLUT_MPORT_737_en = reset;
  assign cosLUT_MPORT_738_data = 32'h3ed95beb;
  assign cosLUT_MPORT_738_addr = 11'h2e2;
  assign cosLUT_MPORT_738_mask = 1'h1;
  assign cosLUT_MPORT_738_en = reset;
  assign cosLUT_MPORT_739_data = 32'h3ed8a5c3;
  assign cosLUT_MPORT_739_addr = 11'h2e3;
  assign cosLUT_MPORT_739_mask = 1'h1;
  assign cosLUT_MPORT_739_en = reset;
  assign cosLUT_MPORT_740_data = 32'h3ed7ef7a;
  assign cosLUT_MPORT_740_addr = 11'h2e4;
  assign cosLUT_MPORT_740_mask = 1'h1;
  assign cosLUT_MPORT_740_en = reset;
  assign cosLUT_MPORT_741_data = 32'h3ed73910;
  assign cosLUT_MPORT_741_addr = 11'h2e5;
  assign cosLUT_MPORT_741_mask = 1'h1;
  assign cosLUT_MPORT_741_en = reset;
  assign cosLUT_MPORT_742_data = 32'h3ed68285;
  assign cosLUT_MPORT_742_addr = 11'h2e6;
  assign cosLUT_MPORT_742_mask = 1'h1;
  assign cosLUT_MPORT_742_en = reset;
  assign cosLUT_MPORT_743_data = 32'h3ed5cbd8;
  assign cosLUT_MPORT_743_addr = 11'h2e7;
  assign cosLUT_MPORT_743_mask = 1'h1;
  assign cosLUT_MPORT_743_en = reset;
  assign cosLUT_MPORT_744_data = 32'h3ed5150b;
  assign cosLUT_MPORT_744_addr = 11'h2e8;
  assign cosLUT_MPORT_744_mask = 1'h1;
  assign cosLUT_MPORT_744_en = reset;
  assign cosLUT_MPORT_745_data = 32'h3ed45e1c;
  assign cosLUT_MPORT_745_addr = 11'h2e9;
  assign cosLUT_MPORT_745_mask = 1'h1;
  assign cosLUT_MPORT_745_en = reset;
  assign cosLUT_MPORT_746_data = 32'h3ed3a70d;
  assign cosLUT_MPORT_746_addr = 11'h2ea;
  assign cosLUT_MPORT_746_mask = 1'h1;
  assign cosLUT_MPORT_746_en = reset;
  assign cosLUT_MPORT_747_data = 32'h3ed2efdd;
  assign cosLUT_MPORT_747_addr = 11'h2eb;
  assign cosLUT_MPORT_747_mask = 1'h1;
  assign cosLUT_MPORT_747_en = reset;
  assign cosLUT_MPORT_748_data = 32'h3ed2388d;
  assign cosLUT_MPORT_748_addr = 11'h2ec;
  assign cosLUT_MPORT_748_mask = 1'h1;
  assign cosLUT_MPORT_748_en = reset;
  assign cosLUT_MPORT_749_data = 32'h3ed1811c;
  assign cosLUT_MPORT_749_addr = 11'h2ed;
  assign cosLUT_MPORT_749_mask = 1'h1;
  assign cosLUT_MPORT_749_en = reset;
  assign cosLUT_MPORT_750_data = 32'h3ed0c98b;
  assign cosLUT_MPORT_750_addr = 11'h2ee;
  assign cosLUT_MPORT_750_mask = 1'h1;
  assign cosLUT_MPORT_750_en = reset;
  assign cosLUT_MPORT_751_data = 32'h3ed011da;
  assign cosLUT_MPORT_751_addr = 11'h2ef;
  assign cosLUT_MPORT_751_mask = 1'h1;
  assign cosLUT_MPORT_751_en = reset;
  assign cosLUT_MPORT_752_data = 32'h3ecf5a08;
  assign cosLUT_MPORT_752_addr = 11'h2f0;
  assign cosLUT_MPORT_752_mask = 1'h1;
  assign cosLUT_MPORT_752_en = reset;
  assign cosLUT_MPORT_753_data = 32'h3ecea217;
  assign cosLUT_MPORT_753_addr = 11'h2f1;
  assign cosLUT_MPORT_753_mask = 1'h1;
  assign cosLUT_MPORT_753_en = reset;
  assign cosLUT_MPORT_754_data = 32'h3ecdea06;
  assign cosLUT_MPORT_754_addr = 11'h2f2;
  assign cosLUT_MPORT_754_mask = 1'h1;
  assign cosLUT_MPORT_754_en = reset;
  assign cosLUT_MPORT_755_data = 32'h3ecd31d4;
  assign cosLUT_MPORT_755_addr = 11'h2f3;
  assign cosLUT_MPORT_755_mask = 1'h1;
  assign cosLUT_MPORT_755_en = reset;
  assign cosLUT_MPORT_756_data = 32'h3ecc7984;
  assign cosLUT_MPORT_756_addr = 11'h2f4;
  assign cosLUT_MPORT_756_mask = 1'h1;
  assign cosLUT_MPORT_756_en = reset;
  assign cosLUT_MPORT_757_data = 32'h3ecbc113;
  assign cosLUT_MPORT_757_addr = 11'h2f5;
  assign cosLUT_MPORT_757_mask = 1'h1;
  assign cosLUT_MPORT_757_en = reset;
  assign cosLUT_MPORT_758_data = 32'h3ecb0884;
  assign cosLUT_MPORT_758_addr = 11'h2f6;
  assign cosLUT_MPORT_758_mask = 1'h1;
  assign cosLUT_MPORT_758_en = reset;
  assign cosLUT_MPORT_759_data = 32'h3eca4fd5;
  assign cosLUT_MPORT_759_addr = 11'h2f7;
  assign cosLUT_MPORT_759_mask = 1'h1;
  assign cosLUT_MPORT_759_en = reset;
  assign cosLUT_MPORT_760_data = 32'h3ec99706;
  assign cosLUT_MPORT_760_addr = 11'h2f8;
  assign cosLUT_MPORT_760_mask = 1'h1;
  assign cosLUT_MPORT_760_en = reset;
  assign cosLUT_MPORT_761_data = 32'h3ec8de19;
  assign cosLUT_MPORT_761_addr = 11'h2f9;
  assign cosLUT_MPORT_761_mask = 1'h1;
  assign cosLUT_MPORT_761_en = reset;
  assign cosLUT_MPORT_762_data = 32'h3ec8250d;
  assign cosLUT_MPORT_762_addr = 11'h2fa;
  assign cosLUT_MPORT_762_mask = 1'h1;
  assign cosLUT_MPORT_762_en = reset;
  assign cosLUT_MPORT_763_data = 32'h3ec76be2;
  assign cosLUT_MPORT_763_addr = 11'h2fb;
  assign cosLUT_MPORT_763_mask = 1'h1;
  assign cosLUT_MPORT_763_en = reset;
  assign cosLUT_MPORT_764_data = 32'h3ec6b298;
  assign cosLUT_MPORT_764_addr = 11'h2fc;
  assign cosLUT_MPORT_764_mask = 1'h1;
  assign cosLUT_MPORT_764_en = reset;
  assign cosLUT_MPORT_765_data = 32'h3ec5f92f;
  assign cosLUT_MPORT_765_addr = 11'h2fd;
  assign cosLUT_MPORT_765_mask = 1'h1;
  assign cosLUT_MPORT_765_en = reset;
  assign cosLUT_MPORT_766_data = 32'h3ec53fa8;
  assign cosLUT_MPORT_766_addr = 11'h2fe;
  assign cosLUT_MPORT_766_mask = 1'h1;
  assign cosLUT_MPORT_766_en = reset;
  assign cosLUT_MPORT_767_data = 32'h3ec48602;
  assign cosLUT_MPORT_767_addr = 11'h2ff;
  assign cosLUT_MPORT_767_mask = 1'h1;
  assign cosLUT_MPORT_767_en = reset;
  assign cosLUT_MPORT_768_data = 32'h3ec3cc3e;
  assign cosLUT_MPORT_768_addr = 11'h300;
  assign cosLUT_MPORT_768_mask = 1'h1;
  assign cosLUT_MPORT_768_en = reset;
  assign cosLUT_MPORT_769_data = 32'h3ec3125c;
  assign cosLUT_MPORT_769_addr = 11'h301;
  assign cosLUT_MPORT_769_mask = 1'h1;
  assign cosLUT_MPORT_769_en = reset;
  assign cosLUT_MPORT_770_data = 32'h3ec2585c;
  assign cosLUT_MPORT_770_addr = 11'h302;
  assign cosLUT_MPORT_770_mask = 1'h1;
  assign cosLUT_MPORT_770_en = reset;
  assign cosLUT_MPORT_771_data = 32'h3ec19e3e;
  assign cosLUT_MPORT_771_addr = 11'h303;
  assign cosLUT_MPORT_771_mask = 1'h1;
  assign cosLUT_MPORT_771_en = reset;
  assign cosLUT_MPORT_772_data = 32'h3ec0e401;
  assign cosLUT_MPORT_772_addr = 11'h304;
  assign cosLUT_MPORT_772_mask = 1'h1;
  assign cosLUT_MPORT_772_en = reset;
  assign cosLUT_MPORT_773_data = 32'h3ec029a8;
  assign cosLUT_MPORT_773_addr = 11'h305;
  assign cosLUT_MPORT_773_mask = 1'h1;
  assign cosLUT_MPORT_773_en = reset;
  assign cosLUT_MPORT_774_data = 32'h3ebf6f30;
  assign cosLUT_MPORT_774_addr = 11'h306;
  assign cosLUT_MPORT_774_mask = 1'h1;
  assign cosLUT_MPORT_774_en = reset;
  assign cosLUT_MPORT_775_data = 32'h3ebeb49b;
  assign cosLUT_MPORT_775_addr = 11'h307;
  assign cosLUT_MPORT_775_mask = 1'h1;
  assign cosLUT_MPORT_775_en = reset;
  assign cosLUT_MPORT_776_data = 32'h3ebdf9e8;
  assign cosLUT_MPORT_776_addr = 11'h308;
  assign cosLUT_MPORT_776_mask = 1'h1;
  assign cosLUT_MPORT_776_en = reset;
  assign cosLUT_MPORT_777_data = 32'h3ebd3f19;
  assign cosLUT_MPORT_777_addr = 11'h309;
  assign cosLUT_MPORT_777_mask = 1'h1;
  assign cosLUT_MPORT_777_en = reset;
  assign cosLUT_MPORT_778_data = 32'h3ebc842c;
  assign cosLUT_MPORT_778_addr = 11'h30a;
  assign cosLUT_MPORT_778_mask = 1'h1;
  assign cosLUT_MPORT_778_en = reset;
  assign cosLUT_MPORT_779_data = 32'h3ebbc922;
  assign cosLUT_MPORT_779_addr = 11'h30b;
  assign cosLUT_MPORT_779_mask = 1'h1;
  assign cosLUT_MPORT_779_en = reset;
  assign cosLUT_MPORT_780_data = 32'h3ebb0dfb;
  assign cosLUT_MPORT_780_addr = 11'h30c;
  assign cosLUT_MPORT_780_mask = 1'h1;
  assign cosLUT_MPORT_780_en = reset;
  assign cosLUT_MPORT_781_data = 32'h3eba52b7;
  assign cosLUT_MPORT_781_addr = 11'h30d;
  assign cosLUT_MPORT_781_mask = 1'h1;
  assign cosLUT_MPORT_781_en = reset;
  assign cosLUT_MPORT_782_data = 32'h3eb99756;
  assign cosLUT_MPORT_782_addr = 11'h30e;
  assign cosLUT_MPORT_782_mask = 1'h1;
  assign cosLUT_MPORT_782_en = reset;
  assign cosLUT_MPORT_783_data = 32'h3eb8dbd9;
  assign cosLUT_MPORT_783_addr = 11'h30f;
  assign cosLUT_MPORT_783_mask = 1'h1;
  assign cosLUT_MPORT_783_en = reset;
  assign cosLUT_MPORT_784_data = 32'h3eb8203f;
  assign cosLUT_MPORT_784_addr = 11'h310;
  assign cosLUT_MPORT_784_mask = 1'h1;
  assign cosLUT_MPORT_784_en = reset;
  assign cosLUT_MPORT_785_data = 32'h3eb76489;
  assign cosLUT_MPORT_785_addr = 11'h311;
  assign cosLUT_MPORT_785_mask = 1'h1;
  assign cosLUT_MPORT_785_en = reset;
  assign cosLUT_MPORT_786_data = 32'h3eb6a8b6;
  assign cosLUT_MPORT_786_addr = 11'h312;
  assign cosLUT_MPORT_786_mask = 1'h1;
  assign cosLUT_MPORT_786_en = reset;
  assign cosLUT_MPORT_787_data = 32'h3eb5ecc7;
  assign cosLUT_MPORT_787_addr = 11'h313;
  assign cosLUT_MPORT_787_mask = 1'h1;
  assign cosLUT_MPORT_787_en = reset;
  assign cosLUT_MPORT_788_data = 32'h3eb530bd;
  assign cosLUT_MPORT_788_addr = 11'h314;
  assign cosLUT_MPORT_788_mask = 1'h1;
  assign cosLUT_MPORT_788_en = reset;
  assign cosLUT_MPORT_789_data = 32'h3eb47496;
  assign cosLUT_MPORT_789_addr = 11'h315;
  assign cosLUT_MPORT_789_mask = 1'h1;
  assign cosLUT_MPORT_789_en = reset;
  assign cosLUT_MPORT_790_data = 32'h3eb3b853;
  assign cosLUT_MPORT_790_addr = 11'h316;
  assign cosLUT_MPORT_790_mask = 1'h1;
  assign cosLUT_MPORT_790_en = reset;
  assign cosLUT_MPORT_791_data = 32'h3eb2fbf5;
  assign cosLUT_MPORT_791_addr = 11'h317;
  assign cosLUT_MPORT_791_mask = 1'h1;
  assign cosLUT_MPORT_791_en = reset;
  assign cosLUT_MPORT_792_data = 32'h3eb23f7b;
  assign cosLUT_MPORT_792_addr = 11'h318;
  assign cosLUT_MPORT_792_mask = 1'h1;
  assign cosLUT_MPORT_792_en = reset;
  assign cosLUT_MPORT_793_data = 32'h3eb182e6;
  assign cosLUT_MPORT_793_addr = 11'h319;
  assign cosLUT_MPORT_793_mask = 1'h1;
  assign cosLUT_MPORT_793_en = reset;
  assign cosLUT_MPORT_794_data = 32'h3eb0c635;
  assign cosLUT_MPORT_794_addr = 11'h31a;
  assign cosLUT_MPORT_794_mask = 1'h1;
  assign cosLUT_MPORT_794_en = reset;
  assign cosLUT_MPORT_795_data = 32'h3eb00969;
  assign cosLUT_MPORT_795_addr = 11'h31b;
  assign cosLUT_MPORT_795_mask = 1'h1;
  assign cosLUT_MPORT_795_en = reset;
  assign cosLUT_MPORT_796_data = 32'h3eaf4c82;
  assign cosLUT_MPORT_796_addr = 11'h31c;
  assign cosLUT_MPORT_796_mask = 1'h1;
  assign cosLUT_MPORT_796_en = reset;
  assign cosLUT_MPORT_797_data = 32'h3eae8f7f;
  assign cosLUT_MPORT_797_addr = 11'h31d;
  assign cosLUT_MPORT_797_mask = 1'h1;
  assign cosLUT_MPORT_797_en = reset;
  assign cosLUT_MPORT_798_data = 32'h3eadd262;
  assign cosLUT_MPORT_798_addr = 11'h31e;
  assign cosLUT_MPORT_798_mask = 1'h1;
  assign cosLUT_MPORT_798_en = reset;
  assign cosLUT_MPORT_799_data = 32'h3ead152a;
  assign cosLUT_MPORT_799_addr = 11'h31f;
  assign cosLUT_MPORT_799_mask = 1'h1;
  assign cosLUT_MPORT_799_en = reset;
  assign cosLUT_MPORT_800_data = 32'h3eac57d7;
  assign cosLUT_MPORT_800_addr = 11'h320;
  assign cosLUT_MPORT_800_mask = 1'h1;
  assign cosLUT_MPORT_800_en = reset;
  assign cosLUT_MPORT_801_data = 32'h3eab9a6a;
  assign cosLUT_MPORT_801_addr = 11'h321;
  assign cosLUT_MPORT_801_mask = 1'h1;
  assign cosLUT_MPORT_801_en = reset;
  assign cosLUT_MPORT_802_data = 32'h3eaadce2;
  assign cosLUT_MPORT_802_addr = 11'h322;
  assign cosLUT_MPORT_802_mask = 1'h1;
  assign cosLUT_MPORT_802_en = reset;
  assign cosLUT_MPORT_803_data = 32'h3eaa1f40;
  assign cosLUT_MPORT_803_addr = 11'h323;
  assign cosLUT_MPORT_803_mask = 1'h1;
  assign cosLUT_MPORT_803_en = reset;
  assign cosLUT_MPORT_804_data = 32'h3ea96184;
  assign cosLUT_MPORT_804_addr = 11'h324;
  assign cosLUT_MPORT_804_mask = 1'h1;
  assign cosLUT_MPORT_804_en = reset;
  assign cosLUT_MPORT_805_data = 32'h3ea8a3ad;
  assign cosLUT_MPORT_805_addr = 11'h325;
  assign cosLUT_MPORT_805_mask = 1'h1;
  assign cosLUT_MPORT_805_en = reset;
  assign cosLUT_MPORT_806_data = 32'h3ea7e5bd;
  assign cosLUT_MPORT_806_addr = 11'h326;
  assign cosLUT_MPORT_806_mask = 1'h1;
  assign cosLUT_MPORT_806_en = reset;
  assign cosLUT_MPORT_807_data = 32'h3ea727b2;
  assign cosLUT_MPORT_807_addr = 11'h327;
  assign cosLUT_MPORT_807_mask = 1'h1;
  assign cosLUT_MPORT_807_en = reset;
  assign cosLUT_MPORT_808_data = 32'h3ea6698e;
  assign cosLUT_MPORT_808_addr = 11'h328;
  assign cosLUT_MPORT_808_mask = 1'h1;
  assign cosLUT_MPORT_808_en = reset;
  assign cosLUT_MPORT_809_data = 32'h3ea5ab50;
  assign cosLUT_MPORT_809_addr = 11'h329;
  assign cosLUT_MPORT_809_mask = 1'h1;
  assign cosLUT_MPORT_809_en = reset;
  assign cosLUT_MPORT_810_data = 32'h3ea4ecf8;
  assign cosLUT_MPORT_810_addr = 11'h32a;
  assign cosLUT_MPORT_810_mask = 1'h1;
  assign cosLUT_MPORT_810_en = reset;
  assign cosLUT_MPORT_811_data = 32'h3ea42e88;
  assign cosLUT_MPORT_811_addr = 11'h32b;
  assign cosLUT_MPORT_811_mask = 1'h1;
  assign cosLUT_MPORT_811_en = reset;
  assign cosLUT_MPORT_812_data = 32'h3ea36ffd;
  assign cosLUT_MPORT_812_addr = 11'h32c;
  assign cosLUT_MPORT_812_mask = 1'h1;
  assign cosLUT_MPORT_812_en = reset;
  assign cosLUT_MPORT_813_data = 32'h3ea2b15a;
  assign cosLUT_MPORT_813_addr = 11'h32d;
  assign cosLUT_MPORT_813_mask = 1'h1;
  assign cosLUT_MPORT_813_en = reset;
  assign cosLUT_MPORT_814_data = 32'h3ea1f29d;
  assign cosLUT_MPORT_814_addr = 11'h32e;
  assign cosLUT_MPORT_814_mask = 1'h1;
  assign cosLUT_MPORT_814_en = reset;
  assign cosLUT_MPORT_815_data = 32'h3ea133c8;
  assign cosLUT_MPORT_815_addr = 11'h32f;
  assign cosLUT_MPORT_815_mask = 1'h1;
  assign cosLUT_MPORT_815_en = reset;
  assign cosLUT_MPORT_816_data = 32'h3ea074d9;
  assign cosLUT_MPORT_816_addr = 11'h330;
  assign cosLUT_MPORT_816_mask = 1'h1;
  assign cosLUT_MPORT_816_en = reset;
  assign cosLUT_MPORT_817_data = 32'h3e9fb5d2;
  assign cosLUT_MPORT_817_addr = 11'h331;
  assign cosLUT_MPORT_817_mask = 1'h1;
  assign cosLUT_MPORT_817_en = reset;
  assign cosLUT_MPORT_818_data = 32'h3e9ef6b2;
  assign cosLUT_MPORT_818_addr = 11'h332;
  assign cosLUT_MPORT_818_mask = 1'h1;
  assign cosLUT_MPORT_818_en = reset;
  assign cosLUT_MPORT_819_data = 32'h3e9e377a;
  assign cosLUT_MPORT_819_addr = 11'h333;
  assign cosLUT_MPORT_819_mask = 1'h1;
  assign cosLUT_MPORT_819_en = reset;
  assign cosLUT_MPORT_820_data = 32'h3e9d7829;
  assign cosLUT_MPORT_820_addr = 11'h334;
  assign cosLUT_MPORT_820_mask = 1'h1;
  assign cosLUT_MPORT_820_en = reset;
  assign cosLUT_MPORT_821_data = 32'h3e9cb8c0;
  assign cosLUT_MPORT_821_addr = 11'h335;
  assign cosLUT_MPORT_821_mask = 1'h1;
  assign cosLUT_MPORT_821_en = reset;
  assign cosLUT_MPORT_822_data = 32'h3e9bf93f;
  assign cosLUT_MPORT_822_addr = 11'h336;
  assign cosLUT_MPORT_822_mask = 1'h1;
  assign cosLUT_MPORT_822_en = reset;
  assign cosLUT_MPORT_823_data = 32'h3e9b39a5;
  assign cosLUT_MPORT_823_addr = 11'h337;
  assign cosLUT_MPORT_823_mask = 1'h1;
  assign cosLUT_MPORT_823_en = reset;
  assign cosLUT_MPORT_824_data = 32'h3e9a79f4;
  assign cosLUT_MPORT_824_addr = 11'h338;
  assign cosLUT_MPORT_824_mask = 1'h1;
  assign cosLUT_MPORT_824_en = reset;
  assign cosLUT_MPORT_825_data = 32'h3e99ba2b;
  assign cosLUT_MPORT_825_addr = 11'h339;
  assign cosLUT_MPORT_825_mask = 1'h1;
  assign cosLUT_MPORT_825_en = reset;
  assign cosLUT_MPORT_826_data = 32'h3e98fa4a;
  assign cosLUT_MPORT_826_addr = 11'h33a;
  assign cosLUT_MPORT_826_mask = 1'h1;
  assign cosLUT_MPORT_826_en = reset;
  assign cosLUT_MPORT_827_data = 32'h3e983a52;
  assign cosLUT_MPORT_827_addr = 11'h33b;
  assign cosLUT_MPORT_827_mask = 1'h1;
  assign cosLUT_MPORT_827_en = reset;
  assign cosLUT_MPORT_828_data = 32'h3e977a42;
  assign cosLUT_MPORT_828_addr = 11'h33c;
  assign cosLUT_MPORT_828_mask = 1'h1;
  assign cosLUT_MPORT_828_en = reset;
  assign cosLUT_MPORT_829_data = 32'h3e96ba1a;
  assign cosLUT_MPORT_829_addr = 11'h33d;
  assign cosLUT_MPORT_829_mask = 1'h1;
  assign cosLUT_MPORT_829_en = reset;
  assign cosLUT_MPORT_830_data = 32'h3e95f9dc;
  assign cosLUT_MPORT_830_addr = 11'h33e;
  assign cosLUT_MPORT_830_mask = 1'h1;
  assign cosLUT_MPORT_830_en = reset;
  assign cosLUT_MPORT_831_data = 32'h3e953986;
  assign cosLUT_MPORT_831_addr = 11'h33f;
  assign cosLUT_MPORT_831_mask = 1'h1;
  assign cosLUT_MPORT_831_en = reset;
  assign cosLUT_MPORT_832_data = 32'h3e94791a;
  assign cosLUT_MPORT_832_addr = 11'h340;
  assign cosLUT_MPORT_832_mask = 1'h1;
  assign cosLUT_MPORT_832_en = reset;
  assign cosLUT_MPORT_833_data = 32'h3e93b896;
  assign cosLUT_MPORT_833_addr = 11'h341;
  assign cosLUT_MPORT_833_mask = 1'h1;
  assign cosLUT_MPORT_833_en = reset;
  assign cosLUT_MPORT_834_data = 32'h3e92f7fc;
  assign cosLUT_MPORT_834_addr = 11'h342;
  assign cosLUT_MPORT_834_mask = 1'h1;
  assign cosLUT_MPORT_834_en = reset;
  assign cosLUT_MPORT_835_data = 32'h3e92374a;
  assign cosLUT_MPORT_835_addr = 11'h343;
  assign cosLUT_MPORT_835_mask = 1'h1;
  assign cosLUT_MPORT_835_en = reset;
  assign cosLUT_MPORT_836_data = 32'h3e917683;
  assign cosLUT_MPORT_836_addr = 11'h344;
  assign cosLUT_MPORT_836_mask = 1'h1;
  assign cosLUT_MPORT_836_en = reset;
  assign cosLUT_MPORT_837_data = 32'h3e90b5a5;
  assign cosLUT_MPORT_837_addr = 11'h345;
  assign cosLUT_MPORT_837_mask = 1'h1;
  assign cosLUT_MPORT_837_en = reset;
  assign cosLUT_MPORT_838_data = 32'h3e8ff4b0;
  assign cosLUT_MPORT_838_addr = 11'h346;
  assign cosLUT_MPORT_838_mask = 1'h1;
  assign cosLUT_MPORT_838_en = reset;
  assign cosLUT_MPORT_839_data = 32'h3e8f33a6;
  assign cosLUT_MPORT_839_addr = 11'h347;
  assign cosLUT_MPORT_839_mask = 1'h1;
  assign cosLUT_MPORT_839_en = reset;
  assign cosLUT_MPORT_840_data = 32'h3e8e7285;
  assign cosLUT_MPORT_840_addr = 11'h348;
  assign cosLUT_MPORT_840_mask = 1'h1;
  assign cosLUT_MPORT_840_en = reset;
  assign cosLUT_MPORT_841_data = 32'h3e8db14e;
  assign cosLUT_MPORT_841_addr = 11'h349;
  assign cosLUT_MPORT_841_mask = 1'h1;
  assign cosLUT_MPORT_841_en = reset;
  assign cosLUT_MPORT_842_data = 32'h3e8cf002;
  assign cosLUT_MPORT_842_addr = 11'h34a;
  assign cosLUT_MPORT_842_mask = 1'h1;
  assign cosLUT_MPORT_842_en = reset;
  assign cosLUT_MPORT_843_data = 32'h3e8c2e9f;
  assign cosLUT_MPORT_843_addr = 11'h34b;
  assign cosLUT_MPORT_843_mask = 1'h1;
  assign cosLUT_MPORT_843_en = reset;
  assign cosLUT_MPORT_844_data = 32'h3e8b6d28;
  assign cosLUT_MPORT_844_addr = 11'h34c;
  assign cosLUT_MPORT_844_mask = 1'h1;
  assign cosLUT_MPORT_844_en = reset;
  assign cosLUT_MPORT_845_data = 32'h3e8aab9a;
  assign cosLUT_MPORT_845_addr = 11'h34d;
  assign cosLUT_MPORT_845_mask = 1'h1;
  assign cosLUT_MPORT_845_en = reset;
  assign cosLUT_MPORT_846_data = 32'h3e89e9f7;
  assign cosLUT_MPORT_846_addr = 11'h34e;
  assign cosLUT_MPORT_846_mask = 1'h1;
  assign cosLUT_MPORT_846_en = reset;
  assign cosLUT_MPORT_847_data = 32'h3e89283f;
  assign cosLUT_MPORT_847_addr = 11'h34f;
  assign cosLUT_MPORT_847_mask = 1'h1;
  assign cosLUT_MPORT_847_en = reset;
  assign cosLUT_MPORT_848_data = 32'h3e886672;
  assign cosLUT_MPORT_848_addr = 11'h350;
  assign cosLUT_MPORT_848_mask = 1'h1;
  assign cosLUT_MPORT_848_en = reset;
  assign cosLUT_MPORT_849_data = 32'h3e87a490;
  assign cosLUT_MPORT_849_addr = 11'h351;
  assign cosLUT_MPORT_849_mask = 1'h1;
  assign cosLUT_MPORT_849_en = reset;
  assign cosLUT_MPORT_850_data = 32'h3e86e298;
  assign cosLUT_MPORT_850_addr = 11'h352;
  assign cosLUT_MPORT_850_mask = 1'h1;
  assign cosLUT_MPORT_850_en = reset;
  assign cosLUT_MPORT_851_data = 32'h3e86208c;
  assign cosLUT_MPORT_851_addr = 11'h353;
  assign cosLUT_MPORT_851_mask = 1'h1;
  assign cosLUT_MPORT_851_en = reset;
  assign cosLUT_MPORT_852_data = 32'h3e855e6b;
  assign cosLUT_MPORT_852_addr = 11'h354;
  assign cosLUT_MPORT_852_mask = 1'h1;
  assign cosLUT_MPORT_852_en = reset;
  assign cosLUT_MPORT_853_data = 32'h3e849c36;
  assign cosLUT_MPORT_853_addr = 11'h355;
  assign cosLUT_MPORT_853_mask = 1'h1;
  assign cosLUT_MPORT_853_en = reset;
  assign cosLUT_MPORT_854_data = 32'h3e83d9ec;
  assign cosLUT_MPORT_854_addr = 11'h356;
  assign cosLUT_MPORT_854_mask = 1'h1;
  assign cosLUT_MPORT_854_en = reset;
  assign cosLUT_MPORT_855_data = 32'h3e83178e;
  assign cosLUT_MPORT_855_addr = 11'h357;
  assign cosLUT_MPORT_855_mask = 1'h1;
  assign cosLUT_MPORT_855_en = reset;
  assign cosLUT_MPORT_856_data = 32'h3e82551c;
  assign cosLUT_MPORT_856_addr = 11'h358;
  assign cosLUT_MPORT_856_mask = 1'h1;
  assign cosLUT_MPORT_856_en = reset;
  assign cosLUT_MPORT_857_data = 32'h3e819295;
  assign cosLUT_MPORT_857_addr = 11'h359;
  assign cosLUT_MPORT_857_mask = 1'h1;
  assign cosLUT_MPORT_857_en = reset;
  assign cosLUT_MPORT_858_data = 32'h3e80cffb;
  assign cosLUT_MPORT_858_addr = 11'h35a;
  assign cosLUT_MPORT_858_mask = 1'h1;
  assign cosLUT_MPORT_858_en = reset;
  assign cosLUT_MPORT_859_data = 32'h3e800d4d;
  assign cosLUT_MPORT_859_addr = 11'h35b;
  assign cosLUT_MPORT_859_mask = 1'h1;
  assign cosLUT_MPORT_859_en = reset;
  assign cosLUT_MPORT_860_data = 32'h3e7e9515;
  assign cosLUT_MPORT_860_addr = 11'h35c;
  assign cosLUT_MPORT_860_mask = 1'h1;
  assign cosLUT_MPORT_860_en = reset;
  assign cosLUT_MPORT_861_data = 32'h3e7d0f6a;
  assign cosLUT_MPORT_861_addr = 11'h35d;
  assign cosLUT_MPORT_861_mask = 1'h1;
  assign cosLUT_MPORT_861_en = reset;
  assign cosLUT_MPORT_862_data = 32'h3e7b8997;
  assign cosLUT_MPORT_862_addr = 11'h35e;
  assign cosLUT_MPORT_862_mask = 1'h1;
  assign cosLUT_MPORT_862_en = reset;
  assign cosLUT_MPORT_863_data = 32'h3e7a039e;
  assign cosLUT_MPORT_863_addr = 11'h35f;
  assign cosLUT_MPORT_863_mask = 1'h1;
  assign cosLUT_MPORT_863_en = reset;
  assign cosLUT_MPORT_864_data = 32'h3e787d7e;
  assign cosLUT_MPORT_864_addr = 11'h360;
  assign cosLUT_MPORT_864_mask = 1'h1;
  assign cosLUT_MPORT_864_en = reset;
  assign cosLUT_MPORT_865_data = 32'h3e76f738;
  assign cosLUT_MPORT_865_addr = 11'h361;
  assign cosLUT_MPORT_865_mask = 1'h1;
  assign cosLUT_MPORT_865_en = reset;
  assign cosLUT_MPORT_866_data = 32'h3e7570cb;
  assign cosLUT_MPORT_866_addr = 11'h362;
  assign cosLUT_MPORT_866_mask = 1'h1;
  assign cosLUT_MPORT_866_en = reset;
  assign cosLUT_MPORT_867_data = 32'h3e73ea39;
  assign cosLUT_MPORT_867_addr = 11'h363;
  assign cosLUT_MPORT_867_mask = 1'h1;
  assign cosLUT_MPORT_867_en = reset;
  assign cosLUT_MPORT_868_data = 32'h3e726381;
  assign cosLUT_MPORT_868_addr = 11'h364;
  assign cosLUT_MPORT_868_mask = 1'h1;
  assign cosLUT_MPORT_868_en = reset;
  assign cosLUT_MPORT_869_data = 32'h3e70dca4;
  assign cosLUT_MPORT_869_addr = 11'h365;
  assign cosLUT_MPORT_869_mask = 1'h1;
  assign cosLUT_MPORT_869_en = reset;
  assign cosLUT_MPORT_870_data = 32'h3e6f55a2;
  assign cosLUT_MPORT_870_addr = 11'h366;
  assign cosLUT_MPORT_870_mask = 1'h1;
  assign cosLUT_MPORT_870_en = reset;
  assign cosLUT_MPORT_871_data = 32'h3e6dce7a;
  assign cosLUT_MPORT_871_addr = 11'h367;
  assign cosLUT_MPORT_871_mask = 1'h1;
  assign cosLUT_MPORT_871_en = reset;
  assign cosLUT_MPORT_872_data = 32'h3e6c472e;
  assign cosLUT_MPORT_872_addr = 11'h368;
  assign cosLUT_MPORT_872_mask = 1'h1;
  assign cosLUT_MPORT_872_en = reset;
  assign cosLUT_MPORT_873_data = 32'h3e6abfbe;
  assign cosLUT_MPORT_873_addr = 11'h369;
  assign cosLUT_MPORT_873_mask = 1'h1;
  assign cosLUT_MPORT_873_en = reset;
  assign cosLUT_MPORT_874_data = 32'h3e693829;
  assign cosLUT_MPORT_874_addr = 11'h36a;
  assign cosLUT_MPORT_874_mask = 1'h1;
  assign cosLUT_MPORT_874_en = reset;
  assign cosLUT_MPORT_875_data = 32'h3e67b071;
  assign cosLUT_MPORT_875_addr = 11'h36b;
  assign cosLUT_MPORT_875_mask = 1'h1;
  assign cosLUT_MPORT_875_en = reset;
  assign cosLUT_MPORT_876_data = 32'h3e662894;
  assign cosLUT_MPORT_876_addr = 11'h36c;
  assign cosLUT_MPORT_876_mask = 1'h1;
  assign cosLUT_MPORT_876_en = reset;
  assign cosLUT_MPORT_877_data = 32'h3e64a094;
  assign cosLUT_MPORT_877_addr = 11'h36d;
  assign cosLUT_MPORT_877_mask = 1'h1;
  assign cosLUT_MPORT_877_en = reset;
  assign cosLUT_MPORT_878_data = 32'h3e631871;
  assign cosLUT_MPORT_878_addr = 11'h36e;
  assign cosLUT_MPORT_878_mask = 1'h1;
  assign cosLUT_MPORT_878_en = reset;
  assign cosLUT_MPORT_879_data = 32'h3e61902b;
  assign cosLUT_MPORT_879_addr = 11'h36f;
  assign cosLUT_MPORT_879_mask = 1'h1;
  assign cosLUT_MPORT_879_en = reset;
  assign cosLUT_MPORT_880_data = 32'h3e6007c2;
  assign cosLUT_MPORT_880_addr = 11'h370;
  assign cosLUT_MPORT_880_mask = 1'h1;
  assign cosLUT_MPORT_880_en = reset;
  assign cosLUT_MPORT_881_data = 32'h3e5e7f36;
  assign cosLUT_MPORT_881_addr = 11'h371;
  assign cosLUT_MPORT_881_mask = 1'h1;
  assign cosLUT_MPORT_881_en = reset;
  assign cosLUT_MPORT_882_data = 32'h3e5cf688;
  assign cosLUT_MPORT_882_addr = 11'h372;
  assign cosLUT_MPORT_882_mask = 1'h1;
  assign cosLUT_MPORT_882_en = reset;
  assign cosLUT_MPORT_883_data = 32'h3e5b6db8;
  assign cosLUT_MPORT_883_addr = 11'h373;
  assign cosLUT_MPORT_883_mask = 1'h1;
  assign cosLUT_MPORT_883_en = reset;
  assign cosLUT_MPORT_884_data = 32'h3e59e4c6;
  assign cosLUT_MPORT_884_addr = 11'h374;
  assign cosLUT_MPORT_884_mask = 1'h1;
  assign cosLUT_MPORT_884_en = reset;
  assign cosLUT_MPORT_885_data = 32'h3e585bb3;
  assign cosLUT_MPORT_885_addr = 11'h375;
  assign cosLUT_MPORT_885_mask = 1'h1;
  assign cosLUT_MPORT_885_en = reset;
  assign cosLUT_MPORT_886_data = 32'h3e56d27e;
  assign cosLUT_MPORT_886_addr = 11'h376;
  assign cosLUT_MPORT_886_mask = 1'h1;
  assign cosLUT_MPORT_886_en = reset;
  assign cosLUT_MPORT_887_data = 32'h3e554928;
  assign cosLUT_MPORT_887_addr = 11'h377;
  assign cosLUT_MPORT_887_mask = 1'h1;
  assign cosLUT_MPORT_887_en = reset;
  assign cosLUT_MPORT_888_data = 32'h3e53bfb1;
  assign cosLUT_MPORT_888_addr = 11'h378;
  assign cosLUT_MPORT_888_mask = 1'h1;
  assign cosLUT_MPORT_888_en = reset;
  assign cosLUT_MPORT_889_data = 32'h3e52361a;
  assign cosLUT_MPORT_889_addr = 11'h379;
  assign cosLUT_MPORT_889_mask = 1'h1;
  assign cosLUT_MPORT_889_en = reset;
  assign cosLUT_MPORT_890_data = 32'h3e50ac61;
  assign cosLUT_MPORT_890_addr = 11'h37a;
  assign cosLUT_MPORT_890_mask = 1'h1;
  assign cosLUT_MPORT_890_en = reset;
  assign cosLUT_MPORT_891_data = 32'h3e4f2289;
  assign cosLUT_MPORT_891_addr = 11'h37b;
  assign cosLUT_MPORT_891_mask = 1'h1;
  assign cosLUT_MPORT_891_en = reset;
  assign cosLUT_MPORT_892_data = 32'h3e4d9891;
  assign cosLUT_MPORT_892_addr = 11'h37c;
  assign cosLUT_MPORT_892_mask = 1'h1;
  assign cosLUT_MPORT_892_en = reset;
  assign cosLUT_MPORT_893_data = 32'h3e4c0e79;
  assign cosLUT_MPORT_893_addr = 11'h37d;
  assign cosLUT_MPORT_893_mask = 1'h1;
  assign cosLUT_MPORT_893_en = reset;
  assign cosLUT_MPORT_894_data = 32'h3e4a8442;
  assign cosLUT_MPORT_894_addr = 11'h37e;
  assign cosLUT_MPORT_894_mask = 1'h1;
  assign cosLUT_MPORT_894_en = reset;
  assign cosLUT_MPORT_895_data = 32'h3e48f9eb;
  assign cosLUT_MPORT_895_addr = 11'h37f;
  assign cosLUT_MPORT_895_mask = 1'h1;
  assign cosLUT_MPORT_895_en = reset;
  assign cosLUT_MPORT_896_data = 32'h3e476f76;
  assign cosLUT_MPORT_896_addr = 11'h380;
  assign cosLUT_MPORT_896_mask = 1'h1;
  assign cosLUT_MPORT_896_en = reset;
  assign cosLUT_MPORT_897_data = 32'h3e45e4e1;
  assign cosLUT_MPORT_897_addr = 11'h381;
  assign cosLUT_MPORT_897_mask = 1'h1;
  assign cosLUT_MPORT_897_en = reset;
  assign cosLUT_MPORT_898_data = 32'h3e445a2e;
  assign cosLUT_MPORT_898_addr = 11'h382;
  assign cosLUT_MPORT_898_mask = 1'h1;
  assign cosLUT_MPORT_898_en = reset;
  assign cosLUT_MPORT_899_data = 32'h3e42cf5d;
  assign cosLUT_MPORT_899_addr = 11'h383;
  assign cosLUT_MPORT_899_mask = 1'h1;
  assign cosLUT_MPORT_899_en = reset;
  assign cosLUT_MPORT_900_data = 32'h3e41446e;
  assign cosLUT_MPORT_900_addr = 11'h384;
  assign cosLUT_MPORT_900_mask = 1'h1;
  assign cosLUT_MPORT_900_en = reset;
  assign cosLUT_MPORT_901_data = 32'h3e3fb961;
  assign cosLUT_MPORT_901_addr = 11'h385;
  assign cosLUT_MPORT_901_mask = 1'h1;
  assign cosLUT_MPORT_901_en = reset;
  assign cosLUT_MPORT_902_data = 32'h3e3e2e36;
  assign cosLUT_MPORT_902_addr = 11'h386;
  assign cosLUT_MPORT_902_mask = 1'h1;
  assign cosLUT_MPORT_902_en = reset;
  assign cosLUT_MPORT_903_data = 32'h3e3ca2ee;
  assign cosLUT_MPORT_903_addr = 11'h387;
  assign cosLUT_MPORT_903_mask = 1'h1;
  assign cosLUT_MPORT_903_en = reset;
  assign cosLUT_MPORT_904_data = 32'h3e3b1789;
  assign cosLUT_MPORT_904_addr = 11'h388;
  assign cosLUT_MPORT_904_mask = 1'h1;
  assign cosLUT_MPORT_904_en = reset;
  assign cosLUT_MPORT_905_data = 32'h3e398c07;
  assign cosLUT_MPORT_905_addr = 11'h389;
  assign cosLUT_MPORT_905_mask = 1'h1;
  assign cosLUT_MPORT_905_en = reset;
  assign cosLUT_MPORT_906_data = 32'h3e380068;
  assign cosLUT_MPORT_906_addr = 11'h38a;
  assign cosLUT_MPORT_906_mask = 1'h1;
  assign cosLUT_MPORT_906_en = reset;
  assign cosLUT_MPORT_907_data = 32'h3e3674ad;
  assign cosLUT_MPORT_907_addr = 11'h38b;
  assign cosLUT_MPORT_907_mask = 1'h1;
  assign cosLUT_MPORT_907_en = reset;
  assign cosLUT_MPORT_908_data = 32'h3e34e8d6;
  assign cosLUT_MPORT_908_addr = 11'h38c;
  assign cosLUT_MPORT_908_mask = 1'h1;
  assign cosLUT_MPORT_908_en = reset;
  assign cosLUT_MPORT_909_data = 32'h3e335ce3;
  assign cosLUT_MPORT_909_addr = 11'h38d;
  assign cosLUT_MPORT_909_mask = 1'h1;
  assign cosLUT_MPORT_909_en = reset;
  assign cosLUT_MPORT_910_data = 32'h3e31d0d4;
  assign cosLUT_MPORT_910_addr = 11'h38e;
  assign cosLUT_MPORT_910_mask = 1'h1;
  assign cosLUT_MPORT_910_en = reset;
  assign cosLUT_MPORT_911_data = 32'h3e3044aa;
  assign cosLUT_MPORT_911_addr = 11'h38f;
  assign cosLUT_MPORT_911_mask = 1'h1;
  assign cosLUT_MPORT_911_en = reset;
  assign cosLUT_MPORT_912_data = 32'h3e2eb864;
  assign cosLUT_MPORT_912_addr = 11'h390;
  assign cosLUT_MPORT_912_mask = 1'h1;
  assign cosLUT_MPORT_912_en = reset;
  assign cosLUT_MPORT_913_data = 32'h3e2d2c04;
  assign cosLUT_MPORT_913_addr = 11'h391;
  assign cosLUT_MPORT_913_mask = 1'h1;
  assign cosLUT_MPORT_913_en = reset;
  assign cosLUT_MPORT_914_data = 32'h3e2b9f89;
  assign cosLUT_MPORT_914_addr = 11'h392;
  assign cosLUT_MPORT_914_mask = 1'h1;
  assign cosLUT_MPORT_914_en = reset;
  assign cosLUT_MPORT_915_data = 32'h3e2a12f3;
  assign cosLUT_MPORT_915_addr = 11'h393;
  assign cosLUT_MPORT_915_mask = 1'h1;
  assign cosLUT_MPORT_915_en = reset;
  assign cosLUT_MPORT_916_data = 32'h3e288644;
  assign cosLUT_MPORT_916_addr = 11'h394;
  assign cosLUT_MPORT_916_mask = 1'h1;
  assign cosLUT_MPORT_916_en = reset;
  assign cosLUT_MPORT_917_data = 32'h3e26f97a;
  assign cosLUT_MPORT_917_addr = 11'h395;
  assign cosLUT_MPORT_917_mask = 1'h1;
  assign cosLUT_MPORT_917_en = reset;
  assign cosLUT_MPORT_918_data = 32'h3e256c96;
  assign cosLUT_MPORT_918_addr = 11'h396;
  assign cosLUT_MPORT_918_mask = 1'h1;
  assign cosLUT_MPORT_918_en = reset;
  assign cosLUT_MPORT_919_data = 32'h3e23df99;
  assign cosLUT_MPORT_919_addr = 11'h397;
  assign cosLUT_MPORT_919_mask = 1'h1;
  assign cosLUT_MPORT_919_en = reset;
  assign cosLUT_MPORT_920_data = 32'h3e225283;
  assign cosLUT_MPORT_920_addr = 11'h398;
  assign cosLUT_MPORT_920_mask = 1'h1;
  assign cosLUT_MPORT_920_en = reset;
  assign cosLUT_MPORT_921_data = 32'h3e20c553;
  assign cosLUT_MPORT_921_addr = 11'h399;
  assign cosLUT_MPORT_921_mask = 1'h1;
  assign cosLUT_MPORT_921_en = reset;
  assign cosLUT_MPORT_922_data = 32'h3e1f380b;
  assign cosLUT_MPORT_922_addr = 11'h39a;
  assign cosLUT_MPORT_922_mask = 1'h1;
  assign cosLUT_MPORT_922_en = reset;
  assign cosLUT_MPORT_923_data = 32'h3e1daaaa;
  assign cosLUT_MPORT_923_addr = 11'h39b;
  assign cosLUT_MPORT_923_mask = 1'h1;
  assign cosLUT_MPORT_923_en = reset;
  assign cosLUT_MPORT_924_data = 32'h3e1c1d31;
  assign cosLUT_MPORT_924_addr = 11'h39c;
  assign cosLUT_MPORT_924_mask = 1'h1;
  assign cosLUT_MPORT_924_en = reset;
  assign cosLUT_MPORT_925_data = 32'h3e1a8fa0;
  assign cosLUT_MPORT_925_addr = 11'h39d;
  assign cosLUT_MPORT_925_mask = 1'h1;
  assign cosLUT_MPORT_925_en = reset;
  assign cosLUT_MPORT_926_data = 32'h3e1901f7;
  assign cosLUT_MPORT_926_addr = 11'h39e;
  assign cosLUT_MPORT_926_mask = 1'h1;
  assign cosLUT_MPORT_926_en = reset;
  assign cosLUT_MPORT_927_data = 32'h3e177436;
  assign cosLUT_MPORT_927_addr = 11'h39f;
  assign cosLUT_MPORT_927_mask = 1'h1;
  assign cosLUT_MPORT_927_en = reset;
  assign cosLUT_MPORT_928_data = 32'h3e15e65e;
  assign cosLUT_MPORT_928_addr = 11'h3a0;
  assign cosLUT_MPORT_928_mask = 1'h1;
  assign cosLUT_MPORT_928_en = reset;
  assign cosLUT_MPORT_929_data = 32'h3e14586f;
  assign cosLUT_MPORT_929_addr = 11'h3a1;
  assign cosLUT_MPORT_929_mask = 1'h1;
  assign cosLUT_MPORT_929_en = reset;
  assign cosLUT_MPORT_930_data = 32'h3e12ca69;
  assign cosLUT_MPORT_930_addr = 11'h3a2;
  assign cosLUT_MPORT_930_mask = 1'h1;
  assign cosLUT_MPORT_930_en = reset;
  assign cosLUT_MPORT_931_data = 32'h3e113c4d;
  assign cosLUT_MPORT_931_addr = 11'h3a3;
  assign cosLUT_MPORT_931_mask = 1'h1;
  assign cosLUT_MPORT_931_en = reset;
  assign cosLUT_MPORT_932_data = 32'h3e0fae1a;
  assign cosLUT_MPORT_932_addr = 11'h3a4;
  assign cosLUT_MPORT_932_mask = 1'h1;
  assign cosLUT_MPORT_932_en = reset;
  assign cosLUT_MPORT_933_data = 32'h3e0e1fd0;
  assign cosLUT_MPORT_933_addr = 11'h3a5;
  assign cosLUT_MPORT_933_mask = 1'h1;
  assign cosLUT_MPORT_933_en = reset;
  assign cosLUT_MPORT_934_data = 32'h3e0c9171;
  assign cosLUT_MPORT_934_addr = 11'h3a6;
  assign cosLUT_MPORT_934_mask = 1'h1;
  assign cosLUT_MPORT_934_en = reset;
  assign cosLUT_MPORT_935_data = 32'h3e0b02fc;
  assign cosLUT_MPORT_935_addr = 11'h3a7;
  assign cosLUT_MPORT_935_mask = 1'h1;
  assign cosLUT_MPORT_935_en = reset;
  assign cosLUT_MPORT_936_data = 32'h3e097472;
  assign cosLUT_MPORT_936_addr = 11'h3a8;
  assign cosLUT_MPORT_936_mask = 1'h1;
  assign cosLUT_MPORT_936_en = reset;
  assign cosLUT_MPORT_937_data = 32'h3e07e5d2;
  assign cosLUT_MPORT_937_addr = 11'h3a9;
  assign cosLUT_MPORT_937_mask = 1'h1;
  assign cosLUT_MPORT_937_en = reset;
  assign cosLUT_MPORT_938_data = 32'h3e06571e;
  assign cosLUT_MPORT_938_addr = 11'h3aa;
  assign cosLUT_MPORT_938_mask = 1'h1;
  assign cosLUT_MPORT_938_en = reset;
  assign cosLUT_MPORT_939_data = 32'h3e04c855;
  assign cosLUT_MPORT_939_addr = 11'h3ab;
  assign cosLUT_MPORT_939_mask = 1'h1;
  assign cosLUT_MPORT_939_en = reset;
  assign cosLUT_MPORT_940_data = 32'h3e033977;
  assign cosLUT_MPORT_940_addr = 11'h3ac;
  assign cosLUT_MPORT_940_mask = 1'h1;
  assign cosLUT_MPORT_940_en = reset;
  assign cosLUT_MPORT_941_data = 32'h3e01aa85;
  assign cosLUT_MPORT_941_addr = 11'h3ad;
  assign cosLUT_MPORT_941_mask = 1'h1;
  assign cosLUT_MPORT_941_en = reset;
  assign cosLUT_MPORT_942_data = 32'h3e001b7f;
  assign cosLUT_MPORT_942_addr = 11'h3ae;
  assign cosLUT_MPORT_942_mask = 1'h1;
  assign cosLUT_MPORT_942_en = reset;
  assign cosLUT_MPORT_943_data = 32'h3dfd18cb;
  assign cosLUT_MPORT_943_addr = 11'h3af;
  assign cosLUT_MPORT_943_mask = 1'h1;
  assign cosLUT_MPORT_943_en = reset;
  assign cosLUT_MPORT_944_data = 32'h3df9fa70;
  assign cosLUT_MPORT_944_addr = 11'h3b0;
  assign cosLUT_MPORT_944_mask = 1'h1;
  assign cosLUT_MPORT_944_en = reset;
  assign cosLUT_MPORT_945_data = 32'h3df6dbef;
  assign cosLUT_MPORT_945_addr = 11'h3b1;
  assign cosLUT_MPORT_945_mask = 1'h1;
  assign cosLUT_MPORT_945_en = reset;
  assign cosLUT_MPORT_946_data = 32'h3df3bd48;
  assign cosLUT_MPORT_946_addr = 11'h3b2;
  assign cosLUT_MPORT_946_mask = 1'h1;
  assign cosLUT_MPORT_946_en = reset;
  assign cosLUT_MPORT_947_data = 32'h3df09e7b;
  assign cosLUT_MPORT_947_addr = 11'h3b3;
  assign cosLUT_MPORT_947_mask = 1'h1;
  assign cosLUT_MPORT_947_en = reset;
  assign cosLUT_MPORT_948_data = 32'h3ded7f8a;
  assign cosLUT_MPORT_948_addr = 11'h3b4;
  assign cosLUT_MPORT_948_mask = 1'h1;
  assign cosLUT_MPORT_948_en = reset;
  assign cosLUT_MPORT_949_data = 32'h3dea6073;
  assign cosLUT_MPORT_949_addr = 11'h3b5;
  assign cosLUT_MPORT_949_mask = 1'h1;
  assign cosLUT_MPORT_949_en = reset;
  assign cosLUT_MPORT_950_data = 32'h3de74138;
  assign cosLUT_MPORT_950_addr = 11'h3b6;
  assign cosLUT_MPORT_950_mask = 1'h1;
  assign cosLUT_MPORT_950_en = reset;
  assign cosLUT_MPORT_951_data = 32'h3de421da;
  assign cosLUT_MPORT_951_addr = 11'h3b7;
  assign cosLUT_MPORT_951_mask = 1'h1;
  assign cosLUT_MPORT_951_en = reset;
  assign cosLUT_MPORT_952_data = 32'h3de10259;
  assign cosLUT_MPORT_952_addr = 11'h3b8;
  assign cosLUT_MPORT_952_mask = 1'h1;
  assign cosLUT_MPORT_952_en = reset;
  assign cosLUT_MPORT_953_data = 32'h3ddde2b4;
  assign cosLUT_MPORT_953_addr = 11'h3b9;
  assign cosLUT_MPORT_953_mask = 1'h1;
  assign cosLUT_MPORT_953_en = reset;
  assign cosLUT_MPORT_954_data = 32'h3ddac2ee;
  assign cosLUT_MPORT_954_addr = 11'h3ba;
  assign cosLUT_MPORT_954_mask = 1'h1;
  assign cosLUT_MPORT_954_en = reset;
  assign cosLUT_MPORT_955_data = 32'h3dd7a305;
  assign cosLUT_MPORT_955_addr = 11'h3bb;
  assign cosLUT_MPORT_955_mask = 1'h1;
  assign cosLUT_MPORT_955_en = reset;
  assign cosLUT_MPORT_956_data = 32'h3dd482fc;
  assign cosLUT_MPORT_956_addr = 11'h3bc;
  assign cosLUT_MPORT_956_mask = 1'h1;
  assign cosLUT_MPORT_956_en = reset;
  assign cosLUT_MPORT_957_data = 32'h3dd162d2;
  assign cosLUT_MPORT_957_addr = 11'h3bd;
  assign cosLUT_MPORT_957_mask = 1'h1;
  assign cosLUT_MPORT_957_en = reset;
  assign cosLUT_MPORT_958_data = 32'h3dce4287;
  assign cosLUT_MPORT_958_addr = 11'h3be;
  assign cosLUT_MPORT_958_mask = 1'h1;
  assign cosLUT_MPORT_958_en = reset;
  assign cosLUT_MPORT_959_data = 32'h3dcb221d;
  assign cosLUT_MPORT_959_addr = 11'h3bf;
  assign cosLUT_MPORT_959_mask = 1'h1;
  assign cosLUT_MPORT_959_en = reset;
  assign cosLUT_MPORT_960_data = 32'h3dc80193;
  assign cosLUT_MPORT_960_addr = 11'h3c0;
  assign cosLUT_MPORT_960_mask = 1'h1;
  assign cosLUT_MPORT_960_en = reset;
  assign cosLUT_MPORT_961_data = 32'h3dc4e0ea;
  assign cosLUT_MPORT_961_addr = 11'h3c1;
  assign cosLUT_MPORT_961_mask = 1'h1;
  assign cosLUT_MPORT_961_en = reset;
  assign cosLUT_MPORT_962_data = 32'h3dc1c023;
  assign cosLUT_MPORT_962_addr = 11'h3c2;
  assign cosLUT_MPORT_962_mask = 1'h1;
  assign cosLUT_MPORT_962_en = reset;
  assign cosLUT_MPORT_963_data = 32'h3dbe9f3e;
  assign cosLUT_MPORT_963_addr = 11'h3c3;
  assign cosLUT_MPORT_963_mask = 1'h1;
  assign cosLUT_MPORT_963_en = reset;
  assign cosLUT_MPORT_964_data = 32'h3dbb7e3c;
  assign cosLUT_MPORT_964_addr = 11'h3c4;
  assign cosLUT_MPORT_964_mask = 1'h1;
  assign cosLUT_MPORT_964_en = reset;
  assign cosLUT_MPORT_965_data = 32'h3db85d1d;
  assign cosLUT_MPORT_965_addr = 11'h3c5;
  assign cosLUT_MPORT_965_mask = 1'h1;
  assign cosLUT_MPORT_965_en = reset;
  assign cosLUT_MPORT_966_data = 32'h3db53be1;
  assign cosLUT_MPORT_966_addr = 11'h3c6;
  assign cosLUT_MPORT_966_mask = 1'h1;
  assign cosLUT_MPORT_966_en = reset;
  assign cosLUT_MPORT_967_data = 32'h3db21a89;
  assign cosLUT_MPORT_967_addr = 11'h3c7;
  assign cosLUT_MPORT_967_mask = 1'h1;
  assign cosLUT_MPORT_967_en = reset;
  assign cosLUT_MPORT_968_data = 32'h3daef916;
  assign cosLUT_MPORT_968_addr = 11'h3c8;
  assign cosLUT_MPORT_968_mask = 1'h1;
  assign cosLUT_MPORT_968_en = reset;
  assign cosLUT_MPORT_969_data = 32'h3dabd788;
  assign cosLUT_MPORT_969_addr = 11'h3c9;
  assign cosLUT_MPORT_969_mask = 1'h1;
  assign cosLUT_MPORT_969_en = reset;
  assign cosLUT_MPORT_970_data = 32'h3da8b5df;
  assign cosLUT_MPORT_970_addr = 11'h3ca;
  assign cosLUT_MPORT_970_mask = 1'h1;
  assign cosLUT_MPORT_970_en = reset;
  assign cosLUT_MPORT_971_data = 32'h3da5941d;
  assign cosLUT_MPORT_971_addr = 11'h3cb;
  assign cosLUT_MPORT_971_mask = 1'h1;
  assign cosLUT_MPORT_971_en = reset;
  assign cosLUT_MPORT_972_data = 32'h3da27240;
  assign cosLUT_MPORT_972_addr = 11'h3cc;
  assign cosLUT_MPORT_972_mask = 1'h1;
  assign cosLUT_MPORT_972_en = reset;
  assign cosLUT_MPORT_973_data = 32'h3d9f504b;
  assign cosLUT_MPORT_973_addr = 11'h3cd;
  assign cosLUT_MPORT_973_mask = 1'h1;
  assign cosLUT_MPORT_973_en = reset;
  assign cosLUT_MPORT_974_data = 32'h3d9c2e3d;
  assign cosLUT_MPORT_974_addr = 11'h3ce;
  assign cosLUT_MPORT_974_mask = 1'h1;
  assign cosLUT_MPORT_974_en = reset;
  assign cosLUT_MPORT_975_data = 32'h3d990c17;
  assign cosLUT_MPORT_975_addr = 11'h3cf;
  assign cosLUT_MPORT_975_mask = 1'h1;
  assign cosLUT_MPORT_975_en = reset;
  assign cosLUT_MPORT_976_data = 32'h3d95e9da;
  assign cosLUT_MPORT_976_addr = 11'h3d0;
  assign cosLUT_MPORT_976_mask = 1'h1;
  assign cosLUT_MPORT_976_en = reset;
  assign cosLUT_MPORT_977_data = 32'h3d92c785;
  assign cosLUT_MPORT_977_addr = 11'h3d1;
  assign cosLUT_MPORT_977_mask = 1'h1;
  assign cosLUT_MPORT_977_en = reset;
  assign cosLUT_MPORT_978_data = 32'h3d8fa51a;
  assign cosLUT_MPORT_978_addr = 11'h3d2;
  assign cosLUT_MPORT_978_mask = 1'h1;
  assign cosLUT_MPORT_978_en = reset;
  assign cosLUT_MPORT_979_data = 32'h3d8c8298;
  assign cosLUT_MPORT_979_addr = 11'h3d3;
  assign cosLUT_MPORT_979_mask = 1'h1;
  assign cosLUT_MPORT_979_en = reset;
  assign cosLUT_MPORT_980_data = 32'h3d896001;
  assign cosLUT_MPORT_980_addr = 11'h3d4;
  assign cosLUT_MPORT_980_mask = 1'h1;
  assign cosLUT_MPORT_980_en = reset;
  assign cosLUT_MPORT_981_data = 32'h3d863d55;
  assign cosLUT_MPORT_981_addr = 11'h3d5;
  assign cosLUT_MPORT_981_mask = 1'h1;
  assign cosLUT_MPORT_981_en = reset;
  assign cosLUT_MPORT_982_data = 32'h3d831a94;
  assign cosLUT_MPORT_982_addr = 11'h3d6;
  assign cosLUT_MPORT_982_mask = 1'h1;
  assign cosLUT_MPORT_982_en = reset;
  assign cosLUT_MPORT_983_data = 32'h3d7fef7c;
  assign cosLUT_MPORT_983_addr = 11'h3d7;
  assign cosLUT_MPORT_983_mask = 1'h1;
  assign cosLUT_MPORT_983_en = reset;
  assign cosLUT_MPORT_984_data = 32'h3d79a9aa;
  assign cosLUT_MPORT_984_addr = 11'h3d8;
  assign cosLUT_MPORT_984_mask = 1'h1;
  assign cosLUT_MPORT_984_en = reset;
  assign cosLUT_MPORT_985_data = 32'h3d7363b2;
  assign cosLUT_MPORT_985_addr = 11'h3d9;
  assign cosLUT_MPORT_985_mask = 1'h1;
  assign cosLUT_MPORT_985_en = reset;
  assign cosLUT_MPORT_986_data = 32'h3d6d1d93;
  assign cosLUT_MPORT_986_addr = 11'h3da;
  assign cosLUT_MPORT_986_mask = 1'h1;
  assign cosLUT_MPORT_986_en = reset;
  assign cosLUT_MPORT_987_data = 32'h3d66d751;
  assign cosLUT_MPORT_987_addr = 11'h3db;
  assign cosLUT_MPORT_987_mask = 1'h1;
  assign cosLUT_MPORT_987_en = reset;
  assign cosLUT_MPORT_988_data = 32'h3d6090ea;
  assign cosLUT_MPORT_988_addr = 11'h3dc;
  assign cosLUT_MPORT_988_mask = 1'h1;
  assign cosLUT_MPORT_988_en = reset;
  assign cosLUT_MPORT_989_data = 32'h3d5a4a61;
  assign cosLUT_MPORT_989_addr = 11'h3dd;
  assign cosLUT_MPORT_989_mask = 1'h1;
  assign cosLUT_MPORT_989_en = reset;
  assign cosLUT_MPORT_990_data = 32'h3d5403b6;
  assign cosLUT_MPORT_990_addr = 11'h3de;
  assign cosLUT_MPORT_990_mask = 1'h1;
  assign cosLUT_MPORT_990_en = reset;
  assign cosLUT_MPORT_991_data = 32'h3d4dbceb;
  assign cosLUT_MPORT_991_addr = 11'h3df;
  assign cosLUT_MPORT_991_mask = 1'h1;
  assign cosLUT_MPORT_991_en = reset;
  assign cosLUT_MPORT_992_data = 32'h3d477600;
  assign cosLUT_MPORT_992_addr = 11'h3e0;
  assign cosLUT_MPORT_992_mask = 1'h1;
  assign cosLUT_MPORT_992_en = reset;
  assign cosLUT_MPORT_993_data = 32'h3d412ef6;
  assign cosLUT_MPORT_993_addr = 11'h3e1;
  assign cosLUT_MPORT_993_mask = 1'h1;
  assign cosLUT_MPORT_993_en = reset;
  assign cosLUT_MPORT_994_data = 32'h3d3ae7ce;
  assign cosLUT_MPORT_994_addr = 11'h3e2;
  assign cosLUT_MPORT_994_mask = 1'h1;
  assign cosLUT_MPORT_994_en = reset;
  assign cosLUT_MPORT_995_data = 32'h3d34a089;
  assign cosLUT_MPORT_995_addr = 11'h3e3;
  assign cosLUT_MPORT_995_mask = 1'h1;
  assign cosLUT_MPORT_995_en = reset;
  assign cosLUT_MPORT_996_data = 32'h3d2e5929;
  assign cosLUT_MPORT_996_addr = 11'h3e4;
  assign cosLUT_MPORT_996_mask = 1'h1;
  assign cosLUT_MPORT_996_en = reset;
  assign cosLUT_MPORT_997_data = 32'h3d2811ad;
  assign cosLUT_MPORT_997_addr = 11'h3e5;
  assign cosLUT_MPORT_997_mask = 1'h1;
  assign cosLUT_MPORT_997_en = reset;
  assign cosLUT_MPORT_998_data = 32'h3d21ca18;
  assign cosLUT_MPORT_998_addr = 11'h3e6;
  assign cosLUT_MPORT_998_mask = 1'h1;
  assign cosLUT_MPORT_998_en = reset;
  assign cosLUT_MPORT_999_data = 32'h3d1b826a;
  assign cosLUT_MPORT_999_addr = 11'h3e7;
  assign cosLUT_MPORT_999_mask = 1'h1;
  assign cosLUT_MPORT_999_en = reset;
  assign cosLUT_MPORT_1000_data = 32'h3d153aa4;
  assign cosLUT_MPORT_1000_addr = 11'h3e8;
  assign cosLUT_MPORT_1000_mask = 1'h1;
  assign cosLUT_MPORT_1000_en = reset;
  assign cosLUT_MPORT_1001_data = 32'h3d0ef2c6;
  assign cosLUT_MPORT_1001_addr = 11'h3e9;
  assign cosLUT_MPORT_1001_mask = 1'h1;
  assign cosLUT_MPORT_1001_en = reset;
  assign cosLUT_MPORT_1002_data = 32'h3d08aad3;
  assign cosLUT_MPORT_1002_addr = 11'h3ea;
  assign cosLUT_MPORT_1002_mask = 1'h1;
  assign cosLUT_MPORT_1002_en = reset;
  assign cosLUT_MPORT_1003_data = 32'h3d0262cb;
  assign cosLUT_MPORT_1003_addr = 11'h3eb;
  assign cosLUT_MPORT_1003_mask = 1'h1;
  assign cosLUT_MPORT_1003_en = reset;
  assign cosLUT_MPORT_1004_data = 32'h3cf8355c;
  assign cosLUT_MPORT_1004_addr = 11'h3ec;
  assign cosLUT_MPORT_1004_mask = 1'h1;
  assign cosLUT_MPORT_1004_en = reset;
  assign cosLUT_MPORT_1005_data = 32'h3ceba4fd;
  assign cosLUT_MPORT_1005_addr = 11'h3ed;
  assign cosLUT_MPORT_1005_mask = 1'h1;
  assign cosLUT_MPORT_1005_en = reset;
  assign cosLUT_MPORT_1006_data = 32'h3cdf1479;
  assign cosLUT_MPORT_1006_addr = 11'h3ee;
  assign cosLUT_MPORT_1006_mask = 1'h1;
  assign cosLUT_MPORT_1006_en = reset;
  assign cosLUT_MPORT_1007_data = 32'h3cd283d3;
  assign cosLUT_MPORT_1007_addr = 11'h3ef;
  assign cosLUT_MPORT_1007_mask = 1'h1;
  assign cosLUT_MPORT_1007_en = reset;
  assign cosLUT_MPORT_1008_data = 32'h3cc5f30c;
  assign cosLUT_MPORT_1008_addr = 11'h3f0;
  assign cosLUT_MPORT_1008_mask = 1'h1;
  assign cosLUT_MPORT_1008_en = reset;
  assign cosLUT_MPORT_1009_data = 32'h3cb96227;
  assign cosLUT_MPORT_1009_addr = 11'h3f1;
  assign cosLUT_MPORT_1009_mask = 1'h1;
  assign cosLUT_MPORT_1009_en = reset;
  assign cosLUT_MPORT_1010_data = 32'h3cacd125;
  assign cosLUT_MPORT_1010_addr = 11'h3f2;
  assign cosLUT_MPORT_1010_mask = 1'h1;
  assign cosLUT_MPORT_1010_en = reset;
  assign cosLUT_MPORT_1011_data = 32'h3ca04008;
  assign cosLUT_MPORT_1011_addr = 11'h3f3;
  assign cosLUT_MPORT_1011_mask = 1'h1;
  assign cosLUT_MPORT_1011_en = reset;
  assign cosLUT_MPORT_1012_data = 32'h3c93aed3;
  assign cosLUT_MPORT_1012_addr = 11'h3f4;
  assign cosLUT_MPORT_1012_mask = 1'h1;
  assign cosLUT_MPORT_1012_en = reset;
  assign cosLUT_MPORT_1013_data = 32'h3c871d87;
  assign cosLUT_MPORT_1013_addr = 11'h3f5;
  assign cosLUT_MPORT_1013_mask = 1'h1;
  assign cosLUT_MPORT_1013_en = reset;
  assign cosLUT_MPORT_1014_data = 32'h3c75184d;
  assign cosLUT_MPORT_1014_addr = 11'h3f6;
  assign cosLUT_MPORT_1014_mask = 1'h1;
  assign cosLUT_MPORT_1014_en = reset;
  assign cosLUT_MPORT_1015_data = 32'h3c5bf566;
  assign cosLUT_MPORT_1015_addr = 11'h3f7;
  assign cosLUT_MPORT_1015_mask = 1'h1;
  assign cosLUT_MPORT_1015_en = reset;
  assign cosLUT_MPORT_1016_data = 32'h3c42d25c;
  assign cosLUT_MPORT_1016_addr = 11'h3f8;
  assign cosLUT_MPORT_1016_mask = 1'h1;
  assign cosLUT_MPORT_1016_en = reset;
  assign cosLUT_MPORT_1017_data = 32'h3c29af35;
  assign cosLUT_MPORT_1017_addr = 11'h3f9;
  assign cosLUT_MPORT_1017_mask = 1'h1;
  assign cosLUT_MPORT_1017_en = reset;
  assign cosLUT_MPORT_1018_data = 32'h3c108bf3;
  assign cosLUT_MPORT_1018_addr = 11'h3fa;
  assign cosLUT_MPORT_1018_mask = 1'h1;
  assign cosLUT_MPORT_1018_en = reset;
  assign cosLUT_MPORT_1019_data = 32'h3beed136;
  assign cosLUT_MPORT_1019_addr = 11'h3fb;
  assign cosLUT_MPORT_1019_mask = 1'h1;
  assign cosLUT_MPORT_1019_en = reset;
  assign cosLUT_MPORT_1020_data = 32'h3bbc8a61;
  assign cosLUT_MPORT_1020_addr = 11'h3fc;
  assign cosLUT_MPORT_1020_mask = 1'h1;
  assign cosLUT_MPORT_1020_en = reset;
  assign cosLUT_MPORT_1021_data = 32'h3b8a4370;
  assign cosLUT_MPORT_1021_addr = 11'h3fd;
  assign cosLUT_MPORT_1021_mask = 1'h1;
  assign cosLUT_MPORT_1021_en = reset;
  assign cosLUT_MPORT_1022_data = 32'h3b2ff8d1;
  assign cosLUT_MPORT_1022_addr = 11'h3fe;
  assign cosLUT_MPORT_1022_mask = 1'h1;
  assign cosLUT_MPORT_1022_en = reset;
  assign cosLUT_MPORT_1023_data = 32'h3a96d54f;
  assign cosLUT_MPORT_1023_addr = 11'h3ff;
  assign cosLUT_MPORT_1023_mask = 1'h1;
  assign cosLUT_MPORT_1023_en = reset;
  assign cosLUT_MPORT_1024_data = 32'h0;
  assign cosLUT_MPORT_1024_addr = 11'h400;
  assign cosLUT_MPORT_1024_mask = 1'h1;
  assign cosLUT_MPORT_1024_en = reset;
  assign io_sinOut_0 = ENReg ? cosLUT_io_sinOut_0_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_1 = ENReg ? cosLUT_io_sinOut_1_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_2 = ENReg ? cosLUT_io_sinOut_2_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_3 = ENReg ? cosLUT_io_sinOut_3_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_4 = ENReg ? cosLUT_io_sinOut_4_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_5 = ENReg ? cosLUT_io_sinOut_5_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_6 = ENReg ? cosLUT_io_sinOut_6_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_sinOut_7 = ENReg ? cosLUT_io_sinOut_7_MPORT_data : 32'h0; // @[LUTbank2.scala 347:32]
  assign io_cosOut_0 = ENReg ? cosLUT_io_cosOut_0_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_1 = ENReg ? cosLUT_io_cosOut_1_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_2 = ENReg ? cosLUT_io_cosOut_2_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_3 = ENReg ? cosLUT_io_cosOut_3_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_4 = ENReg ? cosLUT_io_cosOut_4_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_5 = ENReg ? cosLUT_io_cosOut_5_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_6 = ENReg ? cosLUT_io_cosOut_6_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_cosOut_7 = ENReg ? cosLUT_io_cosOut_7_MPORT_data : 32'h0; // @[LUTbank2.scala 346:32]
  assign io_ENout = ENReg; // @[LUTbank2.scala 343:14]
  assign io_xFWD_0_0 = ENReg ? xFWDReg_0_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_0_1 = ENReg ? xFWDReg_0_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_1_0 = ENReg ? xFWDReg_1_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_1_1 = ENReg ? xFWDReg_1_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_2_0 = ENReg ? xFWDReg_2_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_2_1 = ENReg ? xFWDReg_2_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_3_0 = ENReg ? xFWDReg_3_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_3_1 = ENReg ? xFWDReg_3_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_4_0 = ENReg ? xFWDReg_4_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_4_1 = ENReg ? xFWDReg_4_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_5_0 = ENReg ? xFWDReg_5_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_5_1 = ENReg ? xFWDReg_5_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_6_0 = ENReg ? xFWDReg_6_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_6_1 = ENReg ? xFWDReg_6_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_xFWD_7_0 = ENReg ? xFWDReg_7_0 : 32'h0; // @[LUTbank2.scala 348:32]
  assign io_xFWD_7_1 = ENReg ? xFWDReg_7_1 : 32'h0; // @[LUTbank2.scala 349:32]
  assign io_signFWD_0_0 = ENReg & signReg_0_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_0_1 = ENReg & signReg_0_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_1_0 = ENReg & signReg_1_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_1_1 = ENReg & signReg_1_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_2_0 = ENReg & signReg_2_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_2_1 = ENReg & signReg_2_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_3_0 = ENReg & signReg_3_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_3_1 = ENReg & signReg_3_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_4_0 = ENReg & signReg_4_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_4_1 = ENReg & signReg_4_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_5_0 = ENReg & signReg_5_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_5_1 = ENReg & signReg_5_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_6_0 = ENReg & signReg_6_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_6_1 = ENReg & signReg_6_1; // @[LUTbank2.scala 351:32]
  assign io_signFWD_7_0 = ENReg & signReg_7_0; // @[LUTbank2.scala 350:32]
  assign io_signFWD_7_1 = ENReg & signReg_7_1; // @[LUTbank2.scala 351:32]
  always @(posedge clock) begin
    if (cosLUT_MPORT_en & cosLUT_MPORT_mask) begin
      cosLUT[cosLUT_MPORT_addr] <= cosLUT_MPORT_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1_en & cosLUT_MPORT_1_mask) begin
      cosLUT[cosLUT_MPORT_1_addr] <= cosLUT_MPORT_1_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_2_en & cosLUT_MPORT_2_mask) begin
      cosLUT[cosLUT_MPORT_2_addr] <= cosLUT_MPORT_2_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_3_en & cosLUT_MPORT_3_mask) begin
      cosLUT[cosLUT_MPORT_3_addr] <= cosLUT_MPORT_3_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_4_en & cosLUT_MPORT_4_mask) begin
      cosLUT[cosLUT_MPORT_4_addr] <= cosLUT_MPORT_4_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_5_en & cosLUT_MPORT_5_mask) begin
      cosLUT[cosLUT_MPORT_5_addr] <= cosLUT_MPORT_5_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_6_en & cosLUT_MPORT_6_mask) begin
      cosLUT[cosLUT_MPORT_6_addr] <= cosLUT_MPORT_6_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_7_en & cosLUT_MPORT_7_mask) begin
      cosLUT[cosLUT_MPORT_7_addr] <= cosLUT_MPORT_7_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_8_en & cosLUT_MPORT_8_mask) begin
      cosLUT[cosLUT_MPORT_8_addr] <= cosLUT_MPORT_8_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_9_en & cosLUT_MPORT_9_mask) begin
      cosLUT[cosLUT_MPORT_9_addr] <= cosLUT_MPORT_9_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_10_en & cosLUT_MPORT_10_mask) begin
      cosLUT[cosLUT_MPORT_10_addr] <= cosLUT_MPORT_10_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_11_en & cosLUT_MPORT_11_mask) begin
      cosLUT[cosLUT_MPORT_11_addr] <= cosLUT_MPORT_11_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_12_en & cosLUT_MPORT_12_mask) begin
      cosLUT[cosLUT_MPORT_12_addr] <= cosLUT_MPORT_12_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_13_en & cosLUT_MPORT_13_mask) begin
      cosLUT[cosLUT_MPORT_13_addr] <= cosLUT_MPORT_13_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_14_en & cosLUT_MPORT_14_mask) begin
      cosLUT[cosLUT_MPORT_14_addr] <= cosLUT_MPORT_14_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_15_en & cosLUT_MPORT_15_mask) begin
      cosLUT[cosLUT_MPORT_15_addr] <= cosLUT_MPORT_15_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_16_en & cosLUT_MPORT_16_mask) begin
      cosLUT[cosLUT_MPORT_16_addr] <= cosLUT_MPORT_16_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_17_en & cosLUT_MPORT_17_mask) begin
      cosLUT[cosLUT_MPORT_17_addr] <= cosLUT_MPORT_17_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_18_en & cosLUT_MPORT_18_mask) begin
      cosLUT[cosLUT_MPORT_18_addr] <= cosLUT_MPORT_18_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_19_en & cosLUT_MPORT_19_mask) begin
      cosLUT[cosLUT_MPORT_19_addr] <= cosLUT_MPORT_19_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_20_en & cosLUT_MPORT_20_mask) begin
      cosLUT[cosLUT_MPORT_20_addr] <= cosLUT_MPORT_20_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_21_en & cosLUT_MPORT_21_mask) begin
      cosLUT[cosLUT_MPORT_21_addr] <= cosLUT_MPORT_21_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_22_en & cosLUT_MPORT_22_mask) begin
      cosLUT[cosLUT_MPORT_22_addr] <= cosLUT_MPORT_22_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_23_en & cosLUT_MPORT_23_mask) begin
      cosLUT[cosLUT_MPORT_23_addr] <= cosLUT_MPORT_23_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_24_en & cosLUT_MPORT_24_mask) begin
      cosLUT[cosLUT_MPORT_24_addr] <= cosLUT_MPORT_24_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_25_en & cosLUT_MPORT_25_mask) begin
      cosLUT[cosLUT_MPORT_25_addr] <= cosLUT_MPORT_25_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_26_en & cosLUT_MPORT_26_mask) begin
      cosLUT[cosLUT_MPORT_26_addr] <= cosLUT_MPORT_26_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_27_en & cosLUT_MPORT_27_mask) begin
      cosLUT[cosLUT_MPORT_27_addr] <= cosLUT_MPORT_27_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_28_en & cosLUT_MPORT_28_mask) begin
      cosLUT[cosLUT_MPORT_28_addr] <= cosLUT_MPORT_28_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_29_en & cosLUT_MPORT_29_mask) begin
      cosLUT[cosLUT_MPORT_29_addr] <= cosLUT_MPORT_29_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_30_en & cosLUT_MPORT_30_mask) begin
      cosLUT[cosLUT_MPORT_30_addr] <= cosLUT_MPORT_30_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_31_en & cosLUT_MPORT_31_mask) begin
      cosLUT[cosLUT_MPORT_31_addr] <= cosLUT_MPORT_31_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_32_en & cosLUT_MPORT_32_mask) begin
      cosLUT[cosLUT_MPORT_32_addr] <= cosLUT_MPORT_32_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_33_en & cosLUT_MPORT_33_mask) begin
      cosLUT[cosLUT_MPORT_33_addr] <= cosLUT_MPORT_33_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_34_en & cosLUT_MPORT_34_mask) begin
      cosLUT[cosLUT_MPORT_34_addr] <= cosLUT_MPORT_34_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_35_en & cosLUT_MPORT_35_mask) begin
      cosLUT[cosLUT_MPORT_35_addr] <= cosLUT_MPORT_35_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_36_en & cosLUT_MPORT_36_mask) begin
      cosLUT[cosLUT_MPORT_36_addr] <= cosLUT_MPORT_36_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_37_en & cosLUT_MPORT_37_mask) begin
      cosLUT[cosLUT_MPORT_37_addr] <= cosLUT_MPORT_37_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_38_en & cosLUT_MPORT_38_mask) begin
      cosLUT[cosLUT_MPORT_38_addr] <= cosLUT_MPORT_38_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_39_en & cosLUT_MPORT_39_mask) begin
      cosLUT[cosLUT_MPORT_39_addr] <= cosLUT_MPORT_39_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_40_en & cosLUT_MPORT_40_mask) begin
      cosLUT[cosLUT_MPORT_40_addr] <= cosLUT_MPORT_40_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_41_en & cosLUT_MPORT_41_mask) begin
      cosLUT[cosLUT_MPORT_41_addr] <= cosLUT_MPORT_41_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_42_en & cosLUT_MPORT_42_mask) begin
      cosLUT[cosLUT_MPORT_42_addr] <= cosLUT_MPORT_42_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_43_en & cosLUT_MPORT_43_mask) begin
      cosLUT[cosLUT_MPORT_43_addr] <= cosLUT_MPORT_43_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_44_en & cosLUT_MPORT_44_mask) begin
      cosLUT[cosLUT_MPORT_44_addr] <= cosLUT_MPORT_44_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_45_en & cosLUT_MPORT_45_mask) begin
      cosLUT[cosLUT_MPORT_45_addr] <= cosLUT_MPORT_45_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_46_en & cosLUT_MPORT_46_mask) begin
      cosLUT[cosLUT_MPORT_46_addr] <= cosLUT_MPORT_46_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_47_en & cosLUT_MPORT_47_mask) begin
      cosLUT[cosLUT_MPORT_47_addr] <= cosLUT_MPORT_47_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_48_en & cosLUT_MPORT_48_mask) begin
      cosLUT[cosLUT_MPORT_48_addr] <= cosLUT_MPORT_48_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_49_en & cosLUT_MPORT_49_mask) begin
      cosLUT[cosLUT_MPORT_49_addr] <= cosLUT_MPORT_49_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_50_en & cosLUT_MPORT_50_mask) begin
      cosLUT[cosLUT_MPORT_50_addr] <= cosLUT_MPORT_50_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_51_en & cosLUT_MPORT_51_mask) begin
      cosLUT[cosLUT_MPORT_51_addr] <= cosLUT_MPORT_51_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_52_en & cosLUT_MPORT_52_mask) begin
      cosLUT[cosLUT_MPORT_52_addr] <= cosLUT_MPORT_52_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_53_en & cosLUT_MPORT_53_mask) begin
      cosLUT[cosLUT_MPORT_53_addr] <= cosLUT_MPORT_53_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_54_en & cosLUT_MPORT_54_mask) begin
      cosLUT[cosLUT_MPORT_54_addr] <= cosLUT_MPORT_54_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_55_en & cosLUT_MPORT_55_mask) begin
      cosLUT[cosLUT_MPORT_55_addr] <= cosLUT_MPORT_55_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_56_en & cosLUT_MPORT_56_mask) begin
      cosLUT[cosLUT_MPORT_56_addr] <= cosLUT_MPORT_56_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_57_en & cosLUT_MPORT_57_mask) begin
      cosLUT[cosLUT_MPORT_57_addr] <= cosLUT_MPORT_57_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_58_en & cosLUT_MPORT_58_mask) begin
      cosLUT[cosLUT_MPORT_58_addr] <= cosLUT_MPORT_58_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_59_en & cosLUT_MPORT_59_mask) begin
      cosLUT[cosLUT_MPORT_59_addr] <= cosLUT_MPORT_59_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_60_en & cosLUT_MPORT_60_mask) begin
      cosLUT[cosLUT_MPORT_60_addr] <= cosLUT_MPORT_60_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_61_en & cosLUT_MPORT_61_mask) begin
      cosLUT[cosLUT_MPORT_61_addr] <= cosLUT_MPORT_61_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_62_en & cosLUT_MPORT_62_mask) begin
      cosLUT[cosLUT_MPORT_62_addr] <= cosLUT_MPORT_62_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_63_en & cosLUT_MPORT_63_mask) begin
      cosLUT[cosLUT_MPORT_63_addr] <= cosLUT_MPORT_63_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_64_en & cosLUT_MPORT_64_mask) begin
      cosLUT[cosLUT_MPORT_64_addr] <= cosLUT_MPORT_64_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_65_en & cosLUT_MPORT_65_mask) begin
      cosLUT[cosLUT_MPORT_65_addr] <= cosLUT_MPORT_65_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_66_en & cosLUT_MPORT_66_mask) begin
      cosLUT[cosLUT_MPORT_66_addr] <= cosLUT_MPORT_66_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_67_en & cosLUT_MPORT_67_mask) begin
      cosLUT[cosLUT_MPORT_67_addr] <= cosLUT_MPORT_67_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_68_en & cosLUT_MPORT_68_mask) begin
      cosLUT[cosLUT_MPORT_68_addr] <= cosLUT_MPORT_68_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_69_en & cosLUT_MPORT_69_mask) begin
      cosLUT[cosLUT_MPORT_69_addr] <= cosLUT_MPORT_69_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_70_en & cosLUT_MPORT_70_mask) begin
      cosLUT[cosLUT_MPORT_70_addr] <= cosLUT_MPORT_70_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_71_en & cosLUT_MPORT_71_mask) begin
      cosLUT[cosLUT_MPORT_71_addr] <= cosLUT_MPORT_71_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_72_en & cosLUT_MPORT_72_mask) begin
      cosLUT[cosLUT_MPORT_72_addr] <= cosLUT_MPORT_72_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_73_en & cosLUT_MPORT_73_mask) begin
      cosLUT[cosLUT_MPORT_73_addr] <= cosLUT_MPORT_73_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_74_en & cosLUT_MPORT_74_mask) begin
      cosLUT[cosLUT_MPORT_74_addr] <= cosLUT_MPORT_74_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_75_en & cosLUT_MPORT_75_mask) begin
      cosLUT[cosLUT_MPORT_75_addr] <= cosLUT_MPORT_75_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_76_en & cosLUT_MPORT_76_mask) begin
      cosLUT[cosLUT_MPORT_76_addr] <= cosLUT_MPORT_76_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_77_en & cosLUT_MPORT_77_mask) begin
      cosLUT[cosLUT_MPORT_77_addr] <= cosLUT_MPORT_77_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_78_en & cosLUT_MPORT_78_mask) begin
      cosLUT[cosLUT_MPORT_78_addr] <= cosLUT_MPORT_78_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_79_en & cosLUT_MPORT_79_mask) begin
      cosLUT[cosLUT_MPORT_79_addr] <= cosLUT_MPORT_79_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_80_en & cosLUT_MPORT_80_mask) begin
      cosLUT[cosLUT_MPORT_80_addr] <= cosLUT_MPORT_80_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_81_en & cosLUT_MPORT_81_mask) begin
      cosLUT[cosLUT_MPORT_81_addr] <= cosLUT_MPORT_81_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_82_en & cosLUT_MPORT_82_mask) begin
      cosLUT[cosLUT_MPORT_82_addr] <= cosLUT_MPORT_82_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_83_en & cosLUT_MPORT_83_mask) begin
      cosLUT[cosLUT_MPORT_83_addr] <= cosLUT_MPORT_83_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_84_en & cosLUT_MPORT_84_mask) begin
      cosLUT[cosLUT_MPORT_84_addr] <= cosLUT_MPORT_84_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_85_en & cosLUT_MPORT_85_mask) begin
      cosLUT[cosLUT_MPORT_85_addr] <= cosLUT_MPORT_85_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_86_en & cosLUT_MPORT_86_mask) begin
      cosLUT[cosLUT_MPORT_86_addr] <= cosLUT_MPORT_86_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_87_en & cosLUT_MPORT_87_mask) begin
      cosLUT[cosLUT_MPORT_87_addr] <= cosLUT_MPORT_87_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_88_en & cosLUT_MPORT_88_mask) begin
      cosLUT[cosLUT_MPORT_88_addr] <= cosLUT_MPORT_88_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_89_en & cosLUT_MPORT_89_mask) begin
      cosLUT[cosLUT_MPORT_89_addr] <= cosLUT_MPORT_89_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_90_en & cosLUT_MPORT_90_mask) begin
      cosLUT[cosLUT_MPORT_90_addr] <= cosLUT_MPORT_90_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_91_en & cosLUT_MPORT_91_mask) begin
      cosLUT[cosLUT_MPORT_91_addr] <= cosLUT_MPORT_91_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_92_en & cosLUT_MPORT_92_mask) begin
      cosLUT[cosLUT_MPORT_92_addr] <= cosLUT_MPORT_92_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_93_en & cosLUT_MPORT_93_mask) begin
      cosLUT[cosLUT_MPORT_93_addr] <= cosLUT_MPORT_93_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_94_en & cosLUT_MPORT_94_mask) begin
      cosLUT[cosLUT_MPORT_94_addr] <= cosLUT_MPORT_94_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_95_en & cosLUT_MPORT_95_mask) begin
      cosLUT[cosLUT_MPORT_95_addr] <= cosLUT_MPORT_95_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_96_en & cosLUT_MPORT_96_mask) begin
      cosLUT[cosLUT_MPORT_96_addr] <= cosLUT_MPORT_96_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_97_en & cosLUT_MPORT_97_mask) begin
      cosLUT[cosLUT_MPORT_97_addr] <= cosLUT_MPORT_97_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_98_en & cosLUT_MPORT_98_mask) begin
      cosLUT[cosLUT_MPORT_98_addr] <= cosLUT_MPORT_98_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_99_en & cosLUT_MPORT_99_mask) begin
      cosLUT[cosLUT_MPORT_99_addr] <= cosLUT_MPORT_99_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_100_en & cosLUT_MPORT_100_mask) begin
      cosLUT[cosLUT_MPORT_100_addr] <= cosLUT_MPORT_100_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_101_en & cosLUT_MPORT_101_mask) begin
      cosLUT[cosLUT_MPORT_101_addr] <= cosLUT_MPORT_101_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_102_en & cosLUT_MPORT_102_mask) begin
      cosLUT[cosLUT_MPORT_102_addr] <= cosLUT_MPORT_102_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_103_en & cosLUT_MPORT_103_mask) begin
      cosLUT[cosLUT_MPORT_103_addr] <= cosLUT_MPORT_103_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_104_en & cosLUT_MPORT_104_mask) begin
      cosLUT[cosLUT_MPORT_104_addr] <= cosLUT_MPORT_104_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_105_en & cosLUT_MPORT_105_mask) begin
      cosLUT[cosLUT_MPORT_105_addr] <= cosLUT_MPORT_105_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_106_en & cosLUT_MPORT_106_mask) begin
      cosLUT[cosLUT_MPORT_106_addr] <= cosLUT_MPORT_106_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_107_en & cosLUT_MPORT_107_mask) begin
      cosLUT[cosLUT_MPORT_107_addr] <= cosLUT_MPORT_107_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_108_en & cosLUT_MPORT_108_mask) begin
      cosLUT[cosLUT_MPORT_108_addr] <= cosLUT_MPORT_108_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_109_en & cosLUT_MPORT_109_mask) begin
      cosLUT[cosLUT_MPORT_109_addr] <= cosLUT_MPORT_109_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_110_en & cosLUT_MPORT_110_mask) begin
      cosLUT[cosLUT_MPORT_110_addr] <= cosLUT_MPORT_110_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_111_en & cosLUT_MPORT_111_mask) begin
      cosLUT[cosLUT_MPORT_111_addr] <= cosLUT_MPORT_111_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_112_en & cosLUT_MPORT_112_mask) begin
      cosLUT[cosLUT_MPORT_112_addr] <= cosLUT_MPORT_112_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_113_en & cosLUT_MPORT_113_mask) begin
      cosLUT[cosLUT_MPORT_113_addr] <= cosLUT_MPORT_113_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_114_en & cosLUT_MPORT_114_mask) begin
      cosLUT[cosLUT_MPORT_114_addr] <= cosLUT_MPORT_114_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_115_en & cosLUT_MPORT_115_mask) begin
      cosLUT[cosLUT_MPORT_115_addr] <= cosLUT_MPORT_115_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_116_en & cosLUT_MPORT_116_mask) begin
      cosLUT[cosLUT_MPORT_116_addr] <= cosLUT_MPORT_116_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_117_en & cosLUT_MPORT_117_mask) begin
      cosLUT[cosLUT_MPORT_117_addr] <= cosLUT_MPORT_117_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_118_en & cosLUT_MPORT_118_mask) begin
      cosLUT[cosLUT_MPORT_118_addr] <= cosLUT_MPORT_118_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_119_en & cosLUT_MPORT_119_mask) begin
      cosLUT[cosLUT_MPORT_119_addr] <= cosLUT_MPORT_119_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_120_en & cosLUT_MPORT_120_mask) begin
      cosLUT[cosLUT_MPORT_120_addr] <= cosLUT_MPORT_120_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_121_en & cosLUT_MPORT_121_mask) begin
      cosLUT[cosLUT_MPORT_121_addr] <= cosLUT_MPORT_121_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_122_en & cosLUT_MPORT_122_mask) begin
      cosLUT[cosLUT_MPORT_122_addr] <= cosLUT_MPORT_122_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_123_en & cosLUT_MPORT_123_mask) begin
      cosLUT[cosLUT_MPORT_123_addr] <= cosLUT_MPORT_123_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_124_en & cosLUT_MPORT_124_mask) begin
      cosLUT[cosLUT_MPORT_124_addr] <= cosLUT_MPORT_124_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_125_en & cosLUT_MPORT_125_mask) begin
      cosLUT[cosLUT_MPORT_125_addr] <= cosLUT_MPORT_125_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_126_en & cosLUT_MPORT_126_mask) begin
      cosLUT[cosLUT_MPORT_126_addr] <= cosLUT_MPORT_126_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_127_en & cosLUT_MPORT_127_mask) begin
      cosLUT[cosLUT_MPORT_127_addr] <= cosLUT_MPORT_127_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_128_en & cosLUT_MPORT_128_mask) begin
      cosLUT[cosLUT_MPORT_128_addr] <= cosLUT_MPORT_128_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_129_en & cosLUT_MPORT_129_mask) begin
      cosLUT[cosLUT_MPORT_129_addr] <= cosLUT_MPORT_129_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_130_en & cosLUT_MPORT_130_mask) begin
      cosLUT[cosLUT_MPORT_130_addr] <= cosLUT_MPORT_130_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_131_en & cosLUT_MPORT_131_mask) begin
      cosLUT[cosLUT_MPORT_131_addr] <= cosLUT_MPORT_131_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_132_en & cosLUT_MPORT_132_mask) begin
      cosLUT[cosLUT_MPORT_132_addr] <= cosLUT_MPORT_132_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_133_en & cosLUT_MPORT_133_mask) begin
      cosLUT[cosLUT_MPORT_133_addr] <= cosLUT_MPORT_133_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_134_en & cosLUT_MPORT_134_mask) begin
      cosLUT[cosLUT_MPORT_134_addr] <= cosLUT_MPORT_134_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_135_en & cosLUT_MPORT_135_mask) begin
      cosLUT[cosLUT_MPORT_135_addr] <= cosLUT_MPORT_135_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_136_en & cosLUT_MPORT_136_mask) begin
      cosLUT[cosLUT_MPORT_136_addr] <= cosLUT_MPORT_136_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_137_en & cosLUT_MPORT_137_mask) begin
      cosLUT[cosLUT_MPORT_137_addr] <= cosLUT_MPORT_137_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_138_en & cosLUT_MPORT_138_mask) begin
      cosLUT[cosLUT_MPORT_138_addr] <= cosLUT_MPORT_138_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_139_en & cosLUT_MPORT_139_mask) begin
      cosLUT[cosLUT_MPORT_139_addr] <= cosLUT_MPORT_139_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_140_en & cosLUT_MPORT_140_mask) begin
      cosLUT[cosLUT_MPORT_140_addr] <= cosLUT_MPORT_140_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_141_en & cosLUT_MPORT_141_mask) begin
      cosLUT[cosLUT_MPORT_141_addr] <= cosLUT_MPORT_141_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_142_en & cosLUT_MPORT_142_mask) begin
      cosLUT[cosLUT_MPORT_142_addr] <= cosLUT_MPORT_142_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_143_en & cosLUT_MPORT_143_mask) begin
      cosLUT[cosLUT_MPORT_143_addr] <= cosLUT_MPORT_143_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_144_en & cosLUT_MPORT_144_mask) begin
      cosLUT[cosLUT_MPORT_144_addr] <= cosLUT_MPORT_144_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_145_en & cosLUT_MPORT_145_mask) begin
      cosLUT[cosLUT_MPORT_145_addr] <= cosLUT_MPORT_145_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_146_en & cosLUT_MPORT_146_mask) begin
      cosLUT[cosLUT_MPORT_146_addr] <= cosLUT_MPORT_146_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_147_en & cosLUT_MPORT_147_mask) begin
      cosLUT[cosLUT_MPORT_147_addr] <= cosLUT_MPORT_147_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_148_en & cosLUT_MPORT_148_mask) begin
      cosLUT[cosLUT_MPORT_148_addr] <= cosLUT_MPORT_148_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_149_en & cosLUT_MPORT_149_mask) begin
      cosLUT[cosLUT_MPORT_149_addr] <= cosLUT_MPORT_149_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_150_en & cosLUT_MPORT_150_mask) begin
      cosLUT[cosLUT_MPORT_150_addr] <= cosLUT_MPORT_150_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_151_en & cosLUT_MPORT_151_mask) begin
      cosLUT[cosLUT_MPORT_151_addr] <= cosLUT_MPORT_151_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_152_en & cosLUT_MPORT_152_mask) begin
      cosLUT[cosLUT_MPORT_152_addr] <= cosLUT_MPORT_152_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_153_en & cosLUT_MPORT_153_mask) begin
      cosLUT[cosLUT_MPORT_153_addr] <= cosLUT_MPORT_153_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_154_en & cosLUT_MPORT_154_mask) begin
      cosLUT[cosLUT_MPORT_154_addr] <= cosLUT_MPORT_154_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_155_en & cosLUT_MPORT_155_mask) begin
      cosLUT[cosLUT_MPORT_155_addr] <= cosLUT_MPORT_155_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_156_en & cosLUT_MPORT_156_mask) begin
      cosLUT[cosLUT_MPORT_156_addr] <= cosLUT_MPORT_156_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_157_en & cosLUT_MPORT_157_mask) begin
      cosLUT[cosLUT_MPORT_157_addr] <= cosLUT_MPORT_157_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_158_en & cosLUT_MPORT_158_mask) begin
      cosLUT[cosLUT_MPORT_158_addr] <= cosLUT_MPORT_158_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_159_en & cosLUT_MPORT_159_mask) begin
      cosLUT[cosLUT_MPORT_159_addr] <= cosLUT_MPORT_159_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_160_en & cosLUT_MPORT_160_mask) begin
      cosLUT[cosLUT_MPORT_160_addr] <= cosLUT_MPORT_160_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_161_en & cosLUT_MPORT_161_mask) begin
      cosLUT[cosLUT_MPORT_161_addr] <= cosLUT_MPORT_161_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_162_en & cosLUT_MPORT_162_mask) begin
      cosLUT[cosLUT_MPORT_162_addr] <= cosLUT_MPORT_162_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_163_en & cosLUT_MPORT_163_mask) begin
      cosLUT[cosLUT_MPORT_163_addr] <= cosLUT_MPORT_163_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_164_en & cosLUT_MPORT_164_mask) begin
      cosLUT[cosLUT_MPORT_164_addr] <= cosLUT_MPORT_164_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_165_en & cosLUT_MPORT_165_mask) begin
      cosLUT[cosLUT_MPORT_165_addr] <= cosLUT_MPORT_165_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_166_en & cosLUT_MPORT_166_mask) begin
      cosLUT[cosLUT_MPORT_166_addr] <= cosLUT_MPORT_166_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_167_en & cosLUT_MPORT_167_mask) begin
      cosLUT[cosLUT_MPORT_167_addr] <= cosLUT_MPORT_167_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_168_en & cosLUT_MPORT_168_mask) begin
      cosLUT[cosLUT_MPORT_168_addr] <= cosLUT_MPORT_168_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_169_en & cosLUT_MPORT_169_mask) begin
      cosLUT[cosLUT_MPORT_169_addr] <= cosLUT_MPORT_169_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_170_en & cosLUT_MPORT_170_mask) begin
      cosLUT[cosLUT_MPORT_170_addr] <= cosLUT_MPORT_170_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_171_en & cosLUT_MPORT_171_mask) begin
      cosLUT[cosLUT_MPORT_171_addr] <= cosLUT_MPORT_171_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_172_en & cosLUT_MPORT_172_mask) begin
      cosLUT[cosLUT_MPORT_172_addr] <= cosLUT_MPORT_172_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_173_en & cosLUT_MPORT_173_mask) begin
      cosLUT[cosLUT_MPORT_173_addr] <= cosLUT_MPORT_173_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_174_en & cosLUT_MPORT_174_mask) begin
      cosLUT[cosLUT_MPORT_174_addr] <= cosLUT_MPORT_174_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_175_en & cosLUT_MPORT_175_mask) begin
      cosLUT[cosLUT_MPORT_175_addr] <= cosLUT_MPORT_175_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_176_en & cosLUT_MPORT_176_mask) begin
      cosLUT[cosLUT_MPORT_176_addr] <= cosLUT_MPORT_176_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_177_en & cosLUT_MPORT_177_mask) begin
      cosLUT[cosLUT_MPORT_177_addr] <= cosLUT_MPORT_177_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_178_en & cosLUT_MPORT_178_mask) begin
      cosLUT[cosLUT_MPORT_178_addr] <= cosLUT_MPORT_178_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_179_en & cosLUT_MPORT_179_mask) begin
      cosLUT[cosLUT_MPORT_179_addr] <= cosLUT_MPORT_179_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_180_en & cosLUT_MPORT_180_mask) begin
      cosLUT[cosLUT_MPORT_180_addr] <= cosLUT_MPORT_180_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_181_en & cosLUT_MPORT_181_mask) begin
      cosLUT[cosLUT_MPORT_181_addr] <= cosLUT_MPORT_181_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_182_en & cosLUT_MPORT_182_mask) begin
      cosLUT[cosLUT_MPORT_182_addr] <= cosLUT_MPORT_182_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_183_en & cosLUT_MPORT_183_mask) begin
      cosLUT[cosLUT_MPORT_183_addr] <= cosLUT_MPORT_183_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_184_en & cosLUT_MPORT_184_mask) begin
      cosLUT[cosLUT_MPORT_184_addr] <= cosLUT_MPORT_184_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_185_en & cosLUT_MPORT_185_mask) begin
      cosLUT[cosLUT_MPORT_185_addr] <= cosLUT_MPORT_185_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_186_en & cosLUT_MPORT_186_mask) begin
      cosLUT[cosLUT_MPORT_186_addr] <= cosLUT_MPORT_186_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_187_en & cosLUT_MPORT_187_mask) begin
      cosLUT[cosLUT_MPORT_187_addr] <= cosLUT_MPORT_187_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_188_en & cosLUT_MPORT_188_mask) begin
      cosLUT[cosLUT_MPORT_188_addr] <= cosLUT_MPORT_188_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_189_en & cosLUT_MPORT_189_mask) begin
      cosLUT[cosLUT_MPORT_189_addr] <= cosLUT_MPORT_189_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_190_en & cosLUT_MPORT_190_mask) begin
      cosLUT[cosLUT_MPORT_190_addr] <= cosLUT_MPORT_190_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_191_en & cosLUT_MPORT_191_mask) begin
      cosLUT[cosLUT_MPORT_191_addr] <= cosLUT_MPORT_191_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_192_en & cosLUT_MPORT_192_mask) begin
      cosLUT[cosLUT_MPORT_192_addr] <= cosLUT_MPORT_192_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_193_en & cosLUT_MPORT_193_mask) begin
      cosLUT[cosLUT_MPORT_193_addr] <= cosLUT_MPORT_193_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_194_en & cosLUT_MPORT_194_mask) begin
      cosLUT[cosLUT_MPORT_194_addr] <= cosLUT_MPORT_194_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_195_en & cosLUT_MPORT_195_mask) begin
      cosLUT[cosLUT_MPORT_195_addr] <= cosLUT_MPORT_195_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_196_en & cosLUT_MPORT_196_mask) begin
      cosLUT[cosLUT_MPORT_196_addr] <= cosLUT_MPORT_196_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_197_en & cosLUT_MPORT_197_mask) begin
      cosLUT[cosLUT_MPORT_197_addr] <= cosLUT_MPORT_197_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_198_en & cosLUT_MPORT_198_mask) begin
      cosLUT[cosLUT_MPORT_198_addr] <= cosLUT_MPORT_198_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_199_en & cosLUT_MPORT_199_mask) begin
      cosLUT[cosLUT_MPORT_199_addr] <= cosLUT_MPORT_199_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_200_en & cosLUT_MPORT_200_mask) begin
      cosLUT[cosLUT_MPORT_200_addr] <= cosLUT_MPORT_200_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_201_en & cosLUT_MPORT_201_mask) begin
      cosLUT[cosLUT_MPORT_201_addr] <= cosLUT_MPORT_201_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_202_en & cosLUT_MPORT_202_mask) begin
      cosLUT[cosLUT_MPORT_202_addr] <= cosLUT_MPORT_202_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_203_en & cosLUT_MPORT_203_mask) begin
      cosLUT[cosLUT_MPORT_203_addr] <= cosLUT_MPORT_203_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_204_en & cosLUT_MPORT_204_mask) begin
      cosLUT[cosLUT_MPORT_204_addr] <= cosLUT_MPORT_204_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_205_en & cosLUT_MPORT_205_mask) begin
      cosLUT[cosLUT_MPORT_205_addr] <= cosLUT_MPORT_205_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_206_en & cosLUT_MPORT_206_mask) begin
      cosLUT[cosLUT_MPORT_206_addr] <= cosLUT_MPORT_206_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_207_en & cosLUT_MPORT_207_mask) begin
      cosLUT[cosLUT_MPORT_207_addr] <= cosLUT_MPORT_207_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_208_en & cosLUT_MPORT_208_mask) begin
      cosLUT[cosLUT_MPORT_208_addr] <= cosLUT_MPORT_208_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_209_en & cosLUT_MPORT_209_mask) begin
      cosLUT[cosLUT_MPORT_209_addr] <= cosLUT_MPORT_209_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_210_en & cosLUT_MPORT_210_mask) begin
      cosLUT[cosLUT_MPORT_210_addr] <= cosLUT_MPORT_210_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_211_en & cosLUT_MPORT_211_mask) begin
      cosLUT[cosLUT_MPORT_211_addr] <= cosLUT_MPORT_211_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_212_en & cosLUT_MPORT_212_mask) begin
      cosLUT[cosLUT_MPORT_212_addr] <= cosLUT_MPORT_212_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_213_en & cosLUT_MPORT_213_mask) begin
      cosLUT[cosLUT_MPORT_213_addr] <= cosLUT_MPORT_213_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_214_en & cosLUT_MPORT_214_mask) begin
      cosLUT[cosLUT_MPORT_214_addr] <= cosLUT_MPORT_214_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_215_en & cosLUT_MPORT_215_mask) begin
      cosLUT[cosLUT_MPORT_215_addr] <= cosLUT_MPORT_215_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_216_en & cosLUT_MPORT_216_mask) begin
      cosLUT[cosLUT_MPORT_216_addr] <= cosLUT_MPORT_216_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_217_en & cosLUT_MPORT_217_mask) begin
      cosLUT[cosLUT_MPORT_217_addr] <= cosLUT_MPORT_217_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_218_en & cosLUT_MPORT_218_mask) begin
      cosLUT[cosLUT_MPORT_218_addr] <= cosLUT_MPORT_218_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_219_en & cosLUT_MPORT_219_mask) begin
      cosLUT[cosLUT_MPORT_219_addr] <= cosLUT_MPORT_219_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_220_en & cosLUT_MPORT_220_mask) begin
      cosLUT[cosLUT_MPORT_220_addr] <= cosLUT_MPORT_220_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_221_en & cosLUT_MPORT_221_mask) begin
      cosLUT[cosLUT_MPORT_221_addr] <= cosLUT_MPORT_221_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_222_en & cosLUT_MPORT_222_mask) begin
      cosLUT[cosLUT_MPORT_222_addr] <= cosLUT_MPORT_222_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_223_en & cosLUT_MPORT_223_mask) begin
      cosLUT[cosLUT_MPORT_223_addr] <= cosLUT_MPORT_223_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_224_en & cosLUT_MPORT_224_mask) begin
      cosLUT[cosLUT_MPORT_224_addr] <= cosLUT_MPORT_224_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_225_en & cosLUT_MPORT_225_mask) begin
      cosLUT[cosLUT_MPORT_225_addr] <= cosLUT_MPORT_225_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_226_en & cosLUT_MPORT_226_mask) begin
      cosLUT[cosLUT_MPORT_226_addr] <= cosLUT_MPORT_226_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_227_en & cosLUT_MPORT_227_mask) begin
      cosLUT[cosLUT_MPORT_227_addr] <= cosLUT_MPORT_227_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_228_en & cosLUT_MPORT_228_mask) begin
      cosLUT[cosLUT_MPORT_228_addr] <= cosLUT_MPORT_228_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_229_en & cosLUT_MPORT_229_mask) begin
      cosLUT[cosLUT_MPORT_229_addr] <= cosLUT_MPORT_229_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_230_en & cosLUT_MPORT_230_mask) begin
      cosLUT[cosLUT_MPORT_230_addr] <= cosLUT_MPORT_230_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_231_en & cosLUT_MPORT_231_mask) begin
      cosLUT[cosLUT_MPORT_231_addr] <= cosLUT_MPORT_231_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_232_en & cosLUT_MPORT_232_mask) begin
      cosLUT[cosLUT_MPORT_232_addr] <= cosLUT_MPORT_232_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_233_en & cosLUT_MPORT_233_mask) begin
      cosLUT[cosLUT_MPORT_233_addr] <= cosLUT_MPORT_233_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_234_en & cosLUT_MPORT_234_mask) begin
      cosLUT[cosLUT_MPORT_234_addr] <= cosLUT_MPORT_234_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_235_en & cosLUT_MPORT_235_mask) begin
      cosLUT[cosLUT_MPORT_235_addr] <= cosLUT_MPORT_235_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_236_en & cosLUT_MPORT_236_mask) begin
      cosLUT[cosLUT_MPORT_236_addr] <= cosLUT_MPORT_236_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_237_en & cosLUT_MPORT_237_mask) begin
      cosLUT[cosLUT_MPORT_237_addr] <= cosLUT_MPORT_237_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_238_en & cosLUT_MPORT_238_mask) begin
      cosLUT[cosLUT_MPORT_238_addr] <= cosLUT_MPORT_238_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_239_en & cosLUT_MPORT_239_mask) begin
      cosLUT[cosLUT_MPORT_239_addr] <= cosLUT_MPORT_239_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_240_en & cosLUT_MPORT_240_mask) begin
      cosLUT[cosLUT_MPORT_240_addr] <= cosLUT_MPORT_240_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_241_en & cosLUT_MPORT_241_mask) begin
      cosLUT[cosLUT_MPORT_241_addr] <= cosLUT_MPORT_241_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_242_en & cosLUT_MPORT_242_mask) begin
      cosLUT[cosLUT_MPORT_242_addr] <= cosLUT_MPORT_242_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_243_en & cosLUT_MPORT_243_mask) begin
      cosLUT[cosLUT_MPORT_243_addr] <= cosLUT_MPORT_243_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_244_en & cosLUT_MPORT_244_mask) begin
      cosLUT[cosLUT_MPORT_244_addr] <= cosLUT_MPORT_244_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_245_en & cosLUT_MPORT_245_mask) begin
      cosLUT[cosLUT_MPORT_245_addr] <= cosLUT_MPORT_245_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_246_en & cosLUT_MPORT_246_mask) begin
      cosLUT[cosLUT_MPORT_246_addr] <= cosLUT_MPORT_246_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_247_en & cosLUT_MPORT_247_mask) begin
      cosLUT[cosLUT_MPORT_247_addr] <= cosLUT_MPORT_247_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_248_en & cosLUT_MPORT_248_mask) begin
      cosLUT[cosLUT_MPORT_248_addr] <= cosLUT_MPORT_248_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_249_en & cosLUT_MPORT_249_mask) begin
      cosLUT[cosLUT_MPORT_249_addr] <= cosLUT_MPORT_249_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_250_en & cosLUT_MPORT_250_mask) begin
      cosLUT[cosLUT_MPORT_250_addr] <= cosLUT_MPORT_250_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_251_en & cosLUT_MPORT_251_mask) begin
      cosLUT[cosLUT_MPORT_251_addr] <= cosLUT_MPORT_251_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_252_en & cosLUT_MPORT_252_mask) begin
      cosLUT[cosLUT_MPORT_252_addr] <= cosLUT_MPORT_252_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_253_en & cosLUT_MPORT_253_mask) begin
      cosLUT[cosLUT_MPORT_253_addr] <= cosLUT_MPORT_253_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_254_en & cosLUT_MPORT_254_mask) begin
      cosLUT[cosLUT_MPORT_254_addr] <= cosLUT_MPORT_254_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_255_en & cosLUT_MPORT_255_mask) begin
      cosLUT[cosLUT_MPORT_255_addr] <= cosLUT_MPORT_255_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_256_en & cosLUT_MPORT_256_mask) begin
      cosLUT[cosLUT_MPORT_256_addr] <= cosLUT_MPORT_256_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_257_en & cosLUT_MPORT_257_mask) begin
      cosLUT[cosLUT_MPORT_257_addr] <= cosLUT_MPORT_257_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_258_en & cosLUT_MPORT_258_mask) begin
      cosLUT[cosLUT_MPORT_258_addr] <= cosLUT_MPORT_258_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_259_en & cosLUT_MPORT_259_mask) begin
      cosLUT[cosLUT_MPORT_259_addr] <= cosLUT_MPORT_259_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_260_en & cosLUT_MPORT_260_mask) begin
      cosLUT[cosLUT_MPORT_260_addr] <= cosLUT_MPORT_260_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_261_en & cosLUT_MPORT_261_mask) begin
      cosLUT[cosLUT_MPORT_261_addr] <= cosLUT_MPORT_261_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_262_en & cosLUT_MPORT_262_mask) begin
      cosLUT[cosLUT_MPORT_262_addr] <= cosLUT_MPORT_262_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_263_en & cosLUT_MPORT_263_mask) begin
      cosLUT[cosLUT_MPORT_263_addr] <= cosLUT_MPORT_263_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_264_en & cosLUT_MPORT_264_mask) begin
      cosLUT[cosLUT_MPORT_264_addr] <= cosLUT_MPORT_264_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_265_en & cosLUT_MPORT_265_mask) begin
      cosLUT[cosLUT_MPORT_265_addr] <= cosLUT_MPORT_265_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_266_en & cosLUT_MPORT_266_mask) begin
      cosLUT[cosLUT_MPORT_266_addr] <= cosLUT_MPORT_266_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_267_en & cosLUT_MPORT_267_mask) begin
      cosLUT[cosLUT_MPORT_267_addr] <= cosLUT_MPORT_267_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_268_en & cosLUT_MPORT_268_mask) begin
      cosLUT[cosLUT_MPORT_268_addr] <= cosLUT_MPORT_268_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_269_en & cosLUT_MPORT_269_mask) begin
      cosLUT[cosLUT_MPORT_269_addr] <= cosLUT_MPORT_269_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_270_en & cosLUT_MPORT_270_mask) begin
      cosLUT[cosLUT_MPORT_270_addr] <= cosLUT_MPORT_270_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_271_en & cosLUT_MPORT_271_mask) begin
      cosLUT[cosLUT_MPORT_271_addr] <= cosLUT_MPORT_271_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_272_en & cosLUT_MPORT_272_mask) begin
      cosLUT[cosLUT_MPORT_272_addr] <= cosLUT_MPORT_272_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_273_en & cosLUT_MPORT_273_mask) begin
      cosLUT[cosLUT_MPORT_273_addr] <= cosLUT_MPORT_273_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_274_en & cosLUT_MPORT_274_mask) begin
      cosLUT[cosLUT_MPORT_274_addr] <= cosLUT_MPORT_274_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_275_en & cosLUT_MPORT_275_mask) begin
      cosLUT[cosLUT_MPORT_275_addr] <= cosLUT_MPORT_275_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_276_en & cosLUT_MPORT_276_mask) begin
      cosLUT[cosLUT_MPORT_276_addr] <= cosLUT_MPORT_276_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_277_en & cosLUT_MPORT_277_mask) begin
      cosLUT[cosLUT_MPORT_277_addr] <= cosLUT_MPORT_277_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_278_en & cosLUT_MPORT_278_mask) begin
      cosLUT[cosLUT_MPORT_278_addr] <= cosLUT_MPORT_278_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_279_en & cosLUT_MPORT_279_mask) begin
      cosLUT[cosLUT_MPORT_279_addr] <= cosLUT_MPORT_279_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_280_en & cosLUT_MPORT_280_mask) begin
      cosLUT[cosLUT_MPORT_280_addr] <= cosLUT_MPORT_280_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_281_en & cosLUT_MPORT_281_mask) begin
      cosLUT[cosLUT_MPORT_281_addr] <= cosLUT_MPORT_281_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_282_en & cosLUT_MPORT_282_mask) begin
      cosLUT[cosLUT_MPORT_282_addr] <= cosLUT_MPORT_282_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_283_en & cosLUT_MPORT_283_mask) begin
      cosLUT[cosLUT_MPORT_283_addr] <= cosLUT_MPORT_283_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_284_en & cosLUT_MPORT_284_mask) begin
      cosLUT[cosLUT_MPORT_284_addr] <= cosLUT_MPORT_284_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_285_en & cosLUT_MPORT_285_mask) begin
      cosLUT[cosLUT_MPORT_285_addr] <= cosLUT_MPORT_285_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_286_en & cosLUT_MPORT_286_mask) begin
      cosLUT[cosLUT_MPORT_286_addr] <= cosLUT_MPORT_286_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_287_en & cosLUT_MPORT_287_mask) begin
      cosLUT[cosLUT_MPORT_287_addr] <= cosLUT_MPORT_287_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_288_en & cosLUT_MPORT_288_mask) begin
      cosLUT[cosLUT_MPORT_288_addr] <= cosLUT_MPORT_288_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_289_en & cosLUT_MPORT_289_mask) begin
      cosLUT[cosLUT_MPORT_289_addr] <= cosLUT_MPORT_289_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_290_en & cosLUT_MPORT_290_mask) begin
      cosLUT[cosLUT_MPORT_290_addr] <= cosLUT_MPORT_290_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_291_en & cosLUT_MPORT_291_mask) begin
      cosLUT[cosLUT_MPORT_291_addr] <= cosLUT_MPORT_291_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_292_en & cosLUT_MPORT_292_mask) begin
      cosLUT[cosLUT_MPORT_292_addr] <= cosLUT_MPORT_292_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_293_en & cosLUT_MPORT_293_mask) begin
      cosLUT[cosLUT_MPORT_293_addr] <= cosLUT_MPORT_293_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_294_en & cosLUT_MPORT_294_mask) begin
      cosLUT[cosLUT_MPORT_294_addr] <= cosLUT_MPORT_294_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_295_en & cosLUT_MPORT_295_mask) begin
      cosLUT[cosLUT_MPORT_295_addr] <= cosLUT_MPORT_295_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_296_en & cosLUT_MPORT_296_mask) begin
      cosLUT[cosLUT_MPORT_296_addr] <= cosLUT_MPORT_296_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_297_en & cosLUT_MPORT_297_mask) begin
      cosLUT[cosLUT_MPORT_297_addr] <= cosLUT_MPORT_297_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_298_en & cosLUT_MPORT_298_mask) begin
      cosLUT[cosLUT_MPORT_298_addr] <= cosLUT_MPORT_298_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_299_en & cosLUT_MPORT_299_mask) begin
      cosLUT[cosLUT_MPORT_299_addr] <= cosLUT_MPORT_299_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_300_en & cosLUT_MPORT_300_mask) begin
      cosLUT[cosLUT_MPORT_300_addr] <= cosLUT_MPORT_300_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_301_en & cosLUT_MPORT_301_mask) begin
      cosLUT[cosLUT_MPORT_301_addr] <= cosLUT_MPORT_301_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_302_en & cosLUT_MPORT_302_mask) begin
      cosLUT[cosLUT_MPORT_302_addr] <= cosLUT_MPORT_302_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_303_en & cosLUT_MPORT_303_mask) begin
      cosLUT[cosLUT_MPORT_303_addr] <= cosLUT_MPORT_303_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_304_en & cosLUT_MPORT_304_mask) begin
      cosLUT[cosLUT_MPORT_304_addr] <= cosLUT_MPORT_304_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_305_en & cosLUT_MPORT_305_mask) begin
      cosLUT[cosLUT_MPORT_305_addr] <= cosLUT_MPORT_305_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_306_en & cosLUT_MPORT_306_mask) begin
      cosLUT[cosLUT_MPORT_306_addr] <= cosLUT_MPORT_306_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_307_en & cosLUT_MPORT_307_mask) begin
      cosLUT[cosLUT_MPORT_307_addr] <= cosLUT_MPORT_307_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_308_en & cosLUT_MPORT_308_mask) begin
      cosLUT[cosLUT_MPORT_308_addr] <= cosLUT_MPORT_308_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_309_en & cosLUT_MPORT_309_mask) begin
      cosLUT[cosLUT_MPORT_309_addr] <= cosLUT_MPORT_309_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_310_en & cosLUT_MPORT_310_mask) begin
      cosLUT[cosLUT_MPORT_310_addr] <= cosLUT_MPORT_310_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_311_en & cosLUT_MPORT_311_mask) begin
      cosLUT[cosLUT_MPORT_311_addr] <= cosLUT_MPORT_311_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_312_en & cosLUT_MPORT_312_mask) begin
      cosLUT[cosLUT_MPORT_312_addr] <= cosLUT_MPORT_312_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_313_en & cosLUT_MPORT_313_mask) begin
      cosLUT[cosLUT_MPORT_313_addr] <= cosLUT_MPORT_313_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_314_en & cosLUT_MPORT_314_mask) begin
      cosLUT[cosLUT_MPORT_314_addr] <= cosLUT_MPORT_314_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_315_en & cosLUT_MPORT_315_mask) begin
      cosLUT[cosLUT_MPORT_315_addr] <= cosLUT_MPORT_315_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_316_en & cosLUT_MPORT_316_mask) begin
      cosLUT[cosLUT_MPORT_316_addr] <= cosLUT_MPORT_316_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_317_en & cosLUT_MPORT_317_mask) begin
      cosLUT[cosLUT_MPORT_317_addr] <= cosLUT_MPORT_317_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_318_en & cosLUT_MPORT_318_mask) begin
      cosLUT[cosLUT_MPORT_318_addr] <= cosLUT_MPORT_318_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_319_en & cosLUT_MPORT_319_mask) begin
      cosLUT[cosLUT_MPORT_319_addr] <= cosLUT_MPORT_319_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_320_en & cosLUT_MPORT_320_mask) begin
      cosLUT[cosLUT_MPORT_320_addr] <= cosLUT_MPORT_320_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_321_en & cosLUT_MPORT_321_mask) begin
      cosLUT[cosLUT_MPORT_321_addr] <= cosLUT_MPORT_321_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_322_en & cosLUT_MPORT_322_mask) begin
      cosLUT[cosLUT_MPORT_322_addr] <= cosLUT_MPORT_322_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_323_en & cosLUT_MPORT_323_mask) begin
      cosLUT[cosLUT_MPORT_323_addr] <= cosLUT_MPORT_323_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_324_en & cosLUT_MPORT_324_mask) begin
      cosLUT[cosLUT_MPORT_324_addr] <= cosLUT_MPORT_324_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_325_en & cosLUT_MPORT_325_mask) begin
      cosLUT[cosLUT_MPORT_325_addr] <= cosLUT_MPORT_325_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_326_en & cosLUT_MPORT_326_mask) begin
      cosLUT[cosLUT_MPORT_326_addr] <= cosLUT_MPORT_326_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_327_en & cosLUT_MPORT_327_mask) begin
      cosLUT[cosLUT_MPORT_327_addr] <= cosLUT_MPORT_327_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_328_en & cosLUT_MPORT_328_mask) begin
      cosLUT[cosLUT_MPORT_328_addr] <= cosLUT_MPORT_328_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_329_en & cosLUT_MPORT_329_mask) begin
      cosLUT[cosLUT_MPORT_329_addr] <= cosLUT_MPORT_329_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_330_en & cosLUT_MPORT_330_mask) begin
      cosLUT[cosLUT_MPORT_330_addr] <= cosLUT_MPORT_330_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_331_en & cosLUT_MPORT_331_mask) begin
      cosLUT[cosLUT_MPORT_331_addr] <= cosLUT_MPORT_331_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_332_en & cosLUT_MPORT_332_mask) begin
      cosLUT[cosLUT_MPORT_332_addr] <= cosLUT_MPORT_332_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_333_en & cosLUT_MPORT_333_mask) begin
      cosLUT[cosLUT_MPORT_333_addr] <= cosLUT_MPORT_333_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_334_en & cosLUT_MPORT_334_mask) begin
      cosLUT[cosLUT_MPORT_334_addr] <= cosLUT_MPORT_334_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_335_en & cosLUT_MPORT_335_mask) begin
      cosLUT[cosLUT_MPORT_335_addr] <= cosLUT_MPORT_335_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_336_en & cosLUT_MPORT_336_mask) begin
      cosLUT[cosLUT_MPORT_336_addr] <= cosLUT_MPORT_336_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_337_en & cosLUT_MPORT_337_mask) begin
      cosLUT[cosLUT_MPORT_337_addr] <= cosLUT_MPORT_337_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_338_en & cosLUT_MPORT_338_mask) begin
      cosLUT[cosLUT_MPORT_338_addr] <= cosLUT_MPORT_338_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_339_en & cosLUT_MPORT_339_mask) begin
      cosLUT[cosLUT_MPORT_339_addr] <= cosLUT_MPORT_339_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_340_en & cosLUT_MPORT_340_mask) begin
      cosLUT[cosLUT_MPORT_340_addr] <= cosLUT_MPORT_340_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_341_en & cosLUT_MPORT_341_mask) begin
      cosLUT[cosLUT_MPORT_341_addr] <= cosLUT_MPORT_341_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_342_en & cosLUT_MPORT_342_mask) begin
      cosLUT[cosLUT_MPORT_342_addr] <= cosLUT_MPORT_342_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_343_en & cosLUT_MPORT_343_mask) begin
      cosLUT[cosLUT_MPORT_343_addr] <= cosLUT_MPORT_343_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_344_en & cosLUT_MPORT_344_mask) begin
      cosLUT[cosLUT_MPORT_344_addr] <= cosLUT_MPORT_344_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_345_en & cosLUT_MPORT_345_mask) begin
      cosLUT[cosLUT_MPORT_345_addr] <= cosLUT_MPORT_345_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_346_en & cosLUT_MPORT_346_mask) begin
      cosLUT[cosLUT_MPORT_346_addr] <= cosLUT_MPORT_346_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_347_en & cosLUT_MPORT_347_mask) begin
      cosLUT[cosLUT_MPORT_347_addr] <= cosLUT_MPORT_347_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_348_en & cosLUT_MPORT_348_mask) begin
      cosLUT[cosLUT_MPORT_348_addr] <= cosLUT_MPORT_348_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_349_en & cosLUT_MPORT_349_mask) begin
      cosLUT[cosLUT_MPORT_349_addr] <= cosLUT_MPORT_349_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_350_en & cosLUT_MPORT_350_mask) begin
      cosLUT[cosLUT_MPORT_350_addr] <= cosLUT_MPORT_350_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_351_en & cosLUT_MPORT_351_mask) begin
      cosLUT[cosLUT_MPORT_351_addr] <= cosLUT_MPORT_351_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_352_en & cosLUT_MPORT_352_mask) begin
      cosLUT[cosLUT_MPORT_352_addr] <= cosLUT_MPORT_352_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_353_en & cosLUT_MPORT_353_mask) begin
      cosLUT[cosLUT_MPORT_353_addr] <= cosLUT_MPORT_353_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_354_en & cosLUT_MPORT_354_mask) begin
      cosLUT[cosLUT_MPORT_354_addr] <= cosLUT_MPORT_354_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_355_en & cosLUT_MPORT_355_mask) begin
      cosLUT[cosLUT_MPORT_355_addr] <= cosLUT_MPORT_355_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_356_en & cosLUT_MPORT_356_mask) begin
      cosLUT[cosLUT_MPORT_356_addr] <= cosLUT_MPORT_356_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_357_en & cosLUT_MPORT_357_mask) begin
      cosLUT[cosLUT_MPORT_357_addr] <= cosLUT_MPORT_357_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_358_en & cosLUT_MPORT_358_mask) begin
      cosLUT[cosLUT_MPORT_358_addr] <= cosLUT_MPORT_358_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_359_en & cosLUT_MPORT_359_mask) begin
      cosLUT[cosLUT_MPORT_359_addr] <= cosLUT_MPORT_359_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_360_en & cosLUT_MPORT_360_mask) begin
      cosLUT[cosLUT_MPORT_360_addr] <= cosLUT_MPORT_360_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_361_en & cosLUT_MPORT_361_mask) begin
      cosLUT[cosLUT_MPORT_361_addr] <= cosLUT_MPORT_361_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_362_en & cosLUT_MPORT_362_mask) begin
      cosLUT[cosLUT_MPORT_362_addr] <= cosLUT_MPORT_362_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_363_en & cosLUT_MPORT_363_mask) begin
      cosLUT[cosLUT_MPORT_363_addr] <= cosLUT_MPORT_363_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_364_en & cosLUT_MPORT_364_mask) begin
      cosLUT[cosLUT_MPORT_364_addr] <= cosLUT_MPORT_364_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_365_en & cosLUT_MPORT_365_mask) begin
      cosLUT[cosLUT_MPORT_365_addr] <= cosLUT_MPORT_365_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_366_en & cosLUT_MPORT_366_mask) begin
      cosLUT[cosLUT_MPORT_366_addr] <= cosLUT_MPORT_366_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_367_en & cosLUT_MPORT_367_mask) begin
      cosLUT[cosLUT_MPORT_367_addr] <= cosLUT_MPORT_367_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_368_en & cosLUT_MPORT_368_mask) begin
      cosLUT[cosLUT_MPORT_368_addr] <= cosLUT_MPORT_368_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_369_en & cosLUT_MPORT_369_mask) begin
      cosLUT[cosLUT_MPORT_369_addr] <= cosLUT_MPORT_369_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_370_en & cosLUT_MPORT_370_mask) begin
      cosLUT[cosLUT_MPORT_370_addr] <= cosLUT_MPORT_370_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_371_en & cosLUT_MPORT_371_mask) begin
      cosLUT[cosLUT_MPORT_371_addr] <= cosLUT_MPORT_371_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_372_en & cosLUT_MPORT_372_mask) begin
      cosLUT[cosLUT_MPORT_372_addr] <= cosLUT_MPORT_372_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_373_en & cosLUT_MPORT_373_mask) begin
      cosLUT[cosLUT_MPORT_373_addr] <= cosLUT_MPORT_373_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_374_en & cosLUT_MPORT_374_mask) begin
      cosLUT[cosLUT_MPORT_374_addr] <= cosLUT_MPORT_374_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_375_en & cosLUT_MPORT_375_mask) begin
      cosLUT[cosLUT_MPORT_375_addr] <= cosLUT_MPORT_375_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_376_en & cosLUT_MPORT_376_mask) begin
      cosLUT[cosLUT_MPORT_376_addr] <= cosLUT_MPORT_376_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_377_en & cosLUT_MPORT_377_mask) begin
      cosLUT[cosLUT_MPORT_377_addr] <= cosLUT_MPORT_377_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_378_en & cosLUT_MPORT_378_mask) begin
      cosLUT[cosLUT_MPORT_378_addr] <= cosLUT_MPORT_378_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_379_en & cosLUT_MPORT_379_mask) begin
      cosLUT[cosLUT_MPORT_379_addr] <= cosLUT_MPORT_379_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_380_en & cosLUT_MPORT_380_mask) begin
      cosLUT[cosLUT_MPORT_380_addr] <= cosLUT_MPORT_380_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_381_en & cosLUT_MPORT_381_mask) begin
      cosLUT[cosLUT_MPORT_381_addr] <= cosLUT_MPORT_381_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_382_en & cosLUT_MPORT_382_mask) begin
      cosLUT[cosLUT_MPORT_382_addr] <= cosLUT_MPORT_382_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_383_en & cosLUT_MPORT_383_mask) begin
      cosLUT[cosLUT_MPORT_383_addr] <= cosLUT_MPORT_383_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_384_en & cosLUT_MPORT_384_mask) begin
      cosLUT[cosLUT_MPORT_384_addr] <= cosLUT_MPORT_384_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_385_en & cosLUT_MPORT_385_mask) begin
      cosLUT[cosLUT_MPORT_385_addr] <= cosLUT_MPORT_385_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_386_en & cosLUT_MPORT_386_mask) begin
      cosLUT[cosLUT_MPORT_386_addr] <= cosLUT_MPORT_386_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_387_en & cosLUT_MPORT_387_mask) begin
      cosLUT[cosLUT_MPORT_387_addr] <= cosLUT_MPORT_387_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_388_en & cosLUT_MPORT_388_mask) begin
      cosLUT[cosLUT_MPORT_388_addr] <= cosLUT_MPORT_388_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_389_en & cosLUT_MPORT_389_mask) begin
      cosLUT[cosLUT_MPORT_389_addr] <= cosLUT_MPORT_389_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_390_en & cosLUT_MPORT_390_mask) begin
      cosLUT[cosLUT_MPORT_390_addr] <= cosLUT_MPORT_390_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_391_en & cosLUT_MPORT_391_mask) begin
      cosLUT[cosLUT_MPORT_391_addr] <= cosLUT_MPORT_391_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_392_en & cosLUT_MPORT_392_mask) begin
      cosLUT[cosLUT_MPORT_392_addr] <= cosLUT_MPORT_392_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_393_en & cosLUT_MPORT_393_mask) begin
      cosLUT[cosLUT_MPORT_393_addr] <= cosLUT_MPORT_393_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_394_en & cosLUT_MPORT_394_mask) begin
      cosLUT[cosLUT_MPORT_394_addr] <= cosLUT_MPORT_394_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_395_en & cosLUT_MPORT_395_mask) begin
      cosLUT[cosLUT_MPORT_395_addr] <= cosLUT_MPORT_395_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_396_en & cosLUT_MPORT_396_mask) begin
      cosLUT[cosLUT_MPORT_396_addr] <= cosLUT_MPORT_396_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_397_en & cosLUT_MPORT_397_mask) begin
      cosLUT[cosLUT_MPORT_397_addr] <= cosLUT_MPORT_397_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_398_en & cosLUT_MPORT_398_mask) begin
      cosLUT[cosLUT_MPORT_398_addr] <= cosLUT_MPORT_398_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_399_en & cosLUT_MPORT_399_mask) begin
      cosLUT[cosLUT_MPORT_399_addr] <= cosLUT_MPORT_399_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_400_en & cosLUT_MPORT_400_mask) begin
      cosLUT[cosLUT_MPORT_400_addr] <= cosLUT_MPORT_400_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_401_en & cosLUT_MPORT_401_mask) begin
      cosLUT[cosLUT_MPORT_401_addr] <= cosLUT_MPORT_401_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_402_en & cosLUT_MPORT_402_mask) begin
      cosLUT[cosLUT_MPORT_402_addr] <= cosLUT_MPORT_402_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_403_en & cosLUT_MPORT_403_mask) begin
      cosLUT[cosLUT_MPORT_403_addr] <= cosLUT_MPORT_403_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_404_en & cosLUT_MPORT_404_mask) begin
      cosLUT[cosLUT_MPORT_404_addr] <= cosLUT_MPORT_404_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_405_en & cosLUT_MPORT_405_mask) begin
      cosLUT[cosLUT_MPORT_405_addr] <= cosLUT_MPORT_405_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_406_en & cosLUT_MPORT_406_mask) begin
      cosLUT[cosLUT_MPORT_406_addr] <= cosLUT_MPORT_406_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_407_en & cosLUT_MPORT_407_mask) begin
      cosLUT[cosLUT_MPORT_407_addr] <= cosLUT_MPORT_407_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_408_en & cosLUT_MPORT_408_mask) begin
      cosLUT[cosLUT_MPORT_408_addr] <= cosLUT_MPORT_408_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_409_en & cosLUT_MPORT_409_mask) begin
      cosLUT[cosLUT_MPORT_409_addr] <= cosLUT_MPORT_409_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_410_en & cosLUT_MPORT_410_mask) begin
      cosLUT[cosLUT_MPORT_410_addr] <= cosLUT_MPORT_410_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_411_en & cosLUT_MPORT_411_mask) begin
      cosLUT[cosLUT_MPORT_411_addr] <= cosLUT_MPORT_411_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_412_en & cosLUT_MPORT_412_mask) begin
      cosLUT[cosLUT_MPORT_412_addr] <= cosLUT_MPORT_412_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_413_en & cosLUT_MPORT_413_mask) begin
      cosLUT[cosLUT_MPORT_413_addr] <= cosLUT_MPORT_413_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_414_en & cosLUT_MPORT_414_mask) begin
      cosLUT[cosLUT_MPORT_414_addr] <= cosLUT_MPORT_414_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_415_en & cosLUT_MPORT_415_mask) begin
      cosLUT[cosLUT_MPORT_415_addr] <= cosLUT_MPORT_415_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_416_en & cosLUT_MPORT_416_mask) begin
      cosLUT[cosLUT_MPORT_416_addr] <= cosLUT_MPORT_416_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_417_en & cosLUT_MPORT_417_mask) begin
      cosLUT[cosLUT_MPORT_417_addr] <= cosLUT_MPORT_417_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_418_en & cosLUT_MPORT_418_mask) begin
      cosLUT[cosLUT_MPORT_418_addr] <= cosLUT_MPORT_418_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_419_en & cosLUT_MPORT_419_mask) begin
      cosLUT[cosLUT_MPORT_419_addr] <= cosLUT_MPORT_419_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_420_en & cosLUT_MPORT_420_mask) begin
      cosLUT[cosLUT_MPORT_420_addr] <= cosLUT_MPORT_420_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_421_en & cosLUT_MPORT_421_mask) begin
      cosLUT[cosLUT_MPORT_421_addr] <= cosLUT_MPORT_421_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_422_en & cosLUT_MPORT_422_mask) begin
      cosLUT[cosLUT_MPORT_422_addr] <= cosLUT_MPORT_422_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_423_en & cosLUT_MPORT_423_mask) begin
      cosLUT[cosLUT_MPORT_423_addr] <= cosLUT_MPORT_423_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_424_en & cosLUT_MPORT_424_mask) begin
      cosLUT[cosLUT_MPORT_424_addr] <= cosLUT_MPORT_424_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_425_en & cosLUT_MPORT_425_mask) begin
      cosLUT[cosLUT_MPORT_425_addr] <= cosLUT_MPORT_425_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_426_en & cosLUT_MPORT_426_mask) begin
      cosLUT[cosLUT_MPORT_426_addr] <= cosLUT_MPORT_426_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_427_en & cosLUT_MPORT_427_mask) begin
      cosLUT[cosLUT_MPORT_427_addr] <= cosLUT_MPORT_427_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_428_en & cosLUT_MPORT_428_mask) begin
      cosLUT[cosLUT_MPORT_428_addr] <= cosLUT_MPORT_428_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_429_en & cosLUT_MPORT_429_mask) begin
      cosLUT[cosLUT_MPORT_429_addr] <= cosLUT_MPORT_429_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_430_en & cosLUT_MPORT_430_mask) begin
      cosLUT[cosLUT_MPORT_430_addr] <= cosLUT_MPORT_430_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_431_en & cosLUT_MPORT_431_mask) begin
      cosLUT[cosLUT_MPORT_431_addr] <= cosLUT_MPORT_431_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_432_en & cosLUT_MPORT_432_mask) begin
      cosLUT[cosLUT_MPORT_432_addr] <= cosLUT_MPORT_432_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_433_en & cosLUT_MPORT_433_mask) begin
      cosLUT[cosLUT_MPORT_433_addr] <= cosLUT_MPORT_433_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_434_en & cosLUT_MPORT_434_mask) begin
      cosLUT[cosLUT_MPORT_434_addr] <= cosLUT_MPORT_434_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_435_en & cosLUT_MPORT_435_mask) begin
      cosLUT[cosLUT_MPORT_435_addr] <= cosLUT_MPORT_435_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_436_en & cosLUT_MPORT_436_mask) begin
      cosLUT[cosLUT_MPORT_436_addr] <= cosLUT_MPORT_436_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_437_en & cosLUT_MPORT_437_mask) begin
      cosLUT[cosLUT_MPORT_437_addr] <= cosLUT_MPORT_437_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_438_en & cosLUT_MPORT_438_mask) begin
      cosLUT[cosLUT_MPORT_438_addr] <= cosLUT_MPORT_438_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_439_en & cosLUT_MPORT_439_mask) begin
      cosLUT[cosLUT_MPORT_439_addr] <= cosLUT_MPORT_439_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_440_en & cosLUT_MPORT_440_mask) begin
      cosLUT[cosLUT_MPORT_440_addr] <= cosLUT_MPORT_440_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_441_en & cosLUT_MPORT_441_mask) begin
      cosLUT[cosLUT_MPORT_441_addr] <= cosLUT_MPORT_441_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_442_en & cosLUT_MPORT_442_mask) begin
      cosLUT[cosLUT_MPORT_442_addr] <= cosLUT_MPORT_442_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_443_en & cosLUT_MPORT_443_mask) begin
      cosLUT[cosLUT_MPORT_443_addr] <= cosLUT_MPORT_443_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_444_en & cosLUT_MPORT_444_mask) begin
      cosLUT[cosLUT_MPORT_444_addr] <= cosLUT_MPORT_444_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_445_en & cosLUT_MPORT_445_mask) begin
      cosLUT[cosLUT_MPORT_445_addr] <= cosLUT_MPORT_445_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_446_en & cosLUT_MPORT_446_mask) begin
      cosLUT[cosLUT_MPORT_446_addr] <= cosLUT_MPORT_446_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_447_en & cosLUT_MPORT_447_mask) begin
      cosLUT[cosLUT_MPORT_447_addr] <= cosLUT_MPORT_447_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_448_en & cosLUT_MPORT_448_mask) begin
      cosLUT[cosLUT_MPORT_448_addr] <= cosLUT_MPORT_448_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_449_en & cosLUT_MPORT_449_mask) begin
      cosLUT[cosLUT_MPORT_449_addr] <= cosLUT_MPORT_449_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_450_en & cosLUT_MPORT_450_mask) begin
      cosLUT[cosLUT_MPORT_450_addr] <= cosLUT_MPORT_450_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_451_en & cosLUT_MPORT_451_mask) begin
      cosLUT[cosLUT_MPORT_451_addr] <= cosLUT_MPORT_451_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_452_en & cosLUT_MPORT_452_mask) begin
      cosLUT[cosLUT_MPORT_452_addr] <= cosLUT_MPORT_452_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_453_en & cosLUT_MPORT_453_mask) begin
      cosLUT[cosLUT_MPORT_453_addr] <= cosLUT_MPORT_453_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_454_en & cosLUT_MPORT_454_mask) begin
      cosLUT[cosLUT_MPORT_454_addr] <= cosLUT_MPORT_454_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_455_en & cosLUT_MPORT_455_mask) begin
      cosLUT[cosLUT_MPORT_455_addr] <= cosLUT_MPORT_455_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_456_en & cosLUT_MPORT_456_mask) begin
      cosLUT[cosLUT_MPORT_456_addr] <= cosLUT_MPORT_456_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_457_en & cosLUT_MPORT_457_mask) begin
      cosLUT[cosLUT_MPORT_457_addr] <= cosLUT_MPORT_457_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_458_en & cosLUT_MPORT_458_mask) begin
      cosLUT[cosLUT_MPORT_458_addr] <= cosLUT_MPORT_458_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_459_en & cosLUT_MPORT_459_mask) begin
      cosLUT[cosLUT_MPORT_459_addr] <= cosLUT_MPORT_459_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_460_en & cosLUT_MPORT_460_mask) begin
      cosLUT[cosLUT_MPORT_460_addr] <= cosLUT_MPORT_460_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_461_en & cosLUT_MPORT_461_mask) begin
      cosLUT[cosLUT_MPORT_461_addr] <= cosLUT_MPORT_461_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_462_en & cosLUT_MPORT_462_mask) begin
      cosLUT[cosLUT_MPORT_462_addr] <= cosLUT_MPORT_462_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_463_en & cosLUT_MPORT_463_mask) begin
      cosLUT[cosLUT_MPORT_463_addr] <= cosLUT_MPORT_463_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_464_en & cosLUT_MPORT_464_mask) begin
      cosLUT[cosLUT_MPORT_464_addr] <= cosLUT_MPORT_464_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_465_en & cosLUT_MPORT_465_mask) begin
      cosLUT[cosLUT_MPORT_465_addr] <= cosLUT_MPORT_465_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_466_en & cosLUT_MPORT_466_mask) begin
      cosLUT[cosLUT_MPORT_466_addr] <= cosLUT_MPORT_466_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_467_en & cosLUT_MPORT_467_mask) begin
      cosLUT[cosLUT_MPORT_467_addr] <= cosLUT_MPORT_467_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_468_en & cosLUT_MPORT_468_mask) begin
      cosLUT[cosLUT_MPORT_468_addr] <= cosLUT_MPORT_468_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_469_en & cosLUT_MPORT_469_mask) begin
      cosLUT[cosLUT_MPORT_469_addr] <= cosLUT_MPORT_469_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_470_en & cosLUT_MPORT_470_mask) begin
      cosLUT[cosLUT_MPORT_470_addr] <= cosLUT_MPORT_470_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_471_en & cosLUT_MPORT_471_mask) begin
      cosLUT[cosLUT_MPORT_471_addr] <= cosLUT_MPORT_471_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_472_en & cosLUT_MPORT_472_mask) begin
      cosLUT[cosLUT_MPORT_472_addr] <= cosLUT_MPORT_472_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_473_en & cosLUT_MPORT_473_mask) begin
      cosLUT[cosLUT_MPORT_473_addr] <= cosLUT_MPORT_473_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_474_en & cosLUT_MPORT_474_mask) begin
      cosLUT[cosLUT_MPORT_474_addr] <= cosLUT_MPORT_474_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_475_en & cosLUT_MPORT_475_mask) begin
      cosLUT[cosLUT_MPORT_475_addr] <= cosLUT_MPORT_475_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_476_en & cosLUT_MPORT_476_mask) begin
      cosLUT[cosLUT_MPORT_476_addr] <= cosLUT_MPORT_476_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_477_en & cosLUT_MPORT_477_mask) begin
      cosLUT[cosLUT_MPORT_477_addr] <= cosLUT_MPORT_477_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_478_en & cosLUT_MPORT_478_mask) begin
      cosLUT[cosLUT_MPORT_478_addr] <= cosLUT_MPORT_478_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_479_en & cosLUT_MPORT_479_mask) begin
      cosLUT[cosLUT_MPORT_479_addr] <= cosLUT_MPORT_479_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_480_en & cosLUT_MPORT_480_mask) begin
      cosLUT[cosLUT_MPORT_480_addr] <= cosLUT_MPORT_480_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_481_en & cosLUT_MPORT_481_mask) begin
      cosLUT[cosLUT_MPORT_481_addr] <= cosLUT_MPORT_481_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_482_en & cosLUT_MPORT_482_mask) begin
      cosLUT[cosLUT_MPORT_482_addr] <= cosLUT_MPORT_482_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_483_en & cosLUT_MPORT_483_mask) begin
      cosLUT[cosLUT_MPORT_483_addr] <= cosLUT_MPORT_483_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_484_en & cosLUT_MPORT_484_mask) begin
      cosLUT[cosLUT_MPORT_484_addr] <= cosLUT_MPORT_484_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_485_en & cosLUT_MPORT_485_mask) begin
      cosLUT[cosLUT_MPORT_485_addr] <= cosLUT_MPORT_485_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_486_en & cosLUT_MPORT_486_mask) begin
      cosLUT[cosLUT_MPORT_486_addr] <= cosLUT_MPORT_486_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_487_en & cosLUT_MPORT_487_mask) begin
      cosLUT[cosLUT_MPORT_487_addr] <= cosLUT_MPORT_487_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_488_en & cosLUT_MPORT_488_mask) begin
      cosLUT[cosLUT_MPORT_488_addr] <= cosLUT_MPORT_488_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_489_en & cosLUT_MPORT_489_mask) begin
      cosLUT[cosLUT_MPORT_489_addr] <= cosLUT_MPORT_489_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_490_en & cosLUT_MPORT_490_mask) begin
      cosLUT[cosLUT_MPORT_490_addr] <= cosLUT_MPORT_490_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_491_en & cosLUT_MPORT_491_mask) begin
      cosLUT[cosLUT_MPORT_491_addr] <= cosLUT_MPORT_491_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_492_en & cosLUT_MPORT_492_mask) begin
      cosLUT[cosLUT_MPORT_492_addr] <= cosLUT_MPORT_492_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_493_en & cosLUT_MPORT_493_mask) begin
      cosLUT[cosLUT_MPORT_493_addr] <= cosLUT_MPORT_493_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_494_en & cosLUT_MPORT_494_mask) begin
      cosLUT[cosLUT_MPORT_494_addr] <= cosLUT_MPORT_494_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_495_en & cosLUT_MPORT_495_mask) begin
      cosLUT[cosLUT_MPORT_495_addr] <= cosLUT_MPORT_495_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_496_en & cosLUT_MPORT_496_mask) begin
      cosLUT[cosLUT_MPORT_496_addr] <= cosLUT_MPORT_496_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_497_en & cosLUT_MPORT_497_mask) begin
      cosLUT[cosLUT_MPORT_497_addr] <= cosLUT_MPORT_497_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_498_en & cosLUT_MPORT_498_mask) begin
      cosLUT[cosLUT_MPORT_498_addr] <= cosLUT_MPORT_498_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_499_en & cosLUT_MPORT_499_mask) begin
      cosLUT[cosLUT_MPORT_499_addr] <= cosLUT_MPORT_499_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_500_en & cosLUT_MPORT_500_mask) begin
      cosLUT[cosLUT_MPORT_500_addr] <= cosLUT_MPORT_500_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_501_en & cosLUT_MPORT_501_mask) begin
      cosLUT[cosLUT_MPORT_501_addr] <= cosLUT_MPORT_501_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_502_en & cosLUT_MPORT_502_mask) begin
      cosLUT[cosLUT_MPORT_502_addr] <= cosLUT_MPORT_502_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_503_en & cosLUT_MPORT_503_mask) begin
      cosLUT[cosLUT_MPORT_503_addr] <= cosLUT_MPORT_503_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_504_en & cosLUT_MPORT_504_mask) begin
      cosLUT[cosLUT_MPORT_504_addr] <= cosLUT_MPORT_504_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_505_en & cosLUT_MPORT_505_mask) begin
      cosLUT[cosLUT_MPORT_505_addr] <= cosLUT_MPORT_505_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_506_en & cosLUT_MPORT_506_mask) begin
      cosLUT[cosLUT_MPORT_506_addr] <= cosLUT_MPORT_506_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_507_en & cosLUT_MPORT_507_mask) begin
      cosLUT[cosLUT_MPORT_507_addr] <= cosLUT_MPORT_507_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_508_en & cosLUT_MPORT_508_mask) begin
      cosLUT[cosLUT_MPORT_508_addr] <= cosLUT_MPORT_508_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_509_en & cosLUT_MPORT_509_mask) begin
      cosLUT[cosLUT_MPORT_509_addr] <= cosLUT_MPORT_509_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_510_en & cosLUT_MPORT_510_mask) begin
      cosLUT[cosLUT_MPORT_510_addr] <= cosLUT_MPORT_510_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_511_en & cosLUT_MPORT_511_mask) begin
      cosLUT[cosLUT_MPORT_511_addr] <= cosLUT_MPORT_511_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_512_en & cosLUT_MPORT_512_mask) begin
      cosLUT[cosLUT_MPORT_512_addr] <= cosLUT_MPORT_512_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_513_en & cosLUT_MPORT_513_mask) begin
      cosLUT[cosLUT_MPORT_513_addr] <= cosLUT_MPORT_513_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_514_en & cosLUT_MPORT_514_mask) begin
      cosLUT[cosLUT_MPORT_514_addr] <= cosLUT_MPORT_514_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_515_en & cosLUT_MPORT_515_mask) begin
      cosLUT[cosLUT_MPORT_515_addr] <= cosLUT_MPORT_515_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_516_en & cosLUT_MPORT_516_mask) begin
      cosLUT[cosLUT_MPORT_516_addr] <= cosLUT_MPORT_516_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_517_en & cosLUT_MPORT_517_mask) begin
      cosLUT[cosLUT_MPORT_517_addr] <= cosLUT_MPORT_517_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_518_en & cosLUT_MPORT_518_mask) begin
      cosLUT[cosLUT_MPORT_518_addr] <= cosLUT_MPORT_518_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_519_en & cosLUT_MPORT_519_mask) begin
      cosLUT[cosLUT_MPORT_519_addr] <= cosLUT_MPORT_519_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_520_en & cosLUT_MPORT_520_mask) begin
      cosLUT[cosLUT_MPORT_520_addr] <= cosLUT_MPORT_520_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_521_en & cosLUT_MPORT_521_mask) begin
      cosLUT[cosLUT_MPORT_521_addr] <= cosLUT_MPORT_521_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_522_en & cosLUT_MPORT_522_mask) begin
      cosLUT[cosLUT_MPORT_522_addr] <= cosLUT_MPORT_522_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_523_en & cosLUT_MPORT_523_mask) begin
      cosLUT[cosLUT_MPORT_523_addr] <= cosLUT_MPORT_523_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_524_en & cosLUT_MPORT_524_mask) begin
      cosLUT[cosLUT_MPORT_524_addr] <= cosLUT_MPORT_524_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_525_en & cosLUT_MPORT_525_mask) begin
      cosLUT[cosLUT_MPORT_525_addr] <= cosLUT_MPORT_525_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_526_en & cosLUT_MPORT_526_mask) begin
      cosLUT[cosLUT_MPORT_526_addr] <= cosLUT_MPORT_526_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_527_en & cosLUT_MPORT_527_mask) begin
      cosLUT[cosLUT_MPORT_527_addr] <= cosLUT_MPORT_527_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_528_en & cosLUT_MPORT_528_mask) begin
      cosLUT[cosLUT_MPORT_528_addr] <= cosLUT_MPORT_528_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_529_en & cosLUT_MPORT_529_mask) begin
      cosLUT[cosLUT_MPORT_529_addr] <= cosLUT_MPORT_529_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_530_en & cosLUT_MPORT_530_mask) begin
      cosLUT[cosLUT_MPORT_530_addr] <= cosLUT_MPORT_530_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_531_en & cosLUT_MPORT_531_mask) begin
      cosLUT[cosLUT_MPORT_531_addr] <= cosLUT_MPORT_531_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_532_en & cosLUT_MPORT_532_mask) begin
      cosLUT[cosLUT_MPORT_532_addr] <= cosLUT_MPORT_532_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_533_en & cosLUT_MPORT_533_mask) begin
      cosLUT[cosLUT_MPORT_533_addr] <= cosLUT_MPORT_533_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_534_en & cosLUT_MPORT_534_mask) begin
      cosLUT[cosLUT_MPORT_534_addr] <= cosLUT_MPORT_534_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_535_en & cosLUT_MPORT_535_mask) begin
      cosLUT[cosLUT_MPORT_535_addr] <= cosLUT_MPORT_535_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_536_en & cosLUT_MPORT_536_mask) begin
      cosLUT[cosLUT_MPORT_536_addr] <= cosLUT_MPORT_536_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_537_en & cosLUT_MPORT_537_mask) begin
      cosLUT[cosLUT_MPORT_537_addr] <= cosLUT_MPORT_537_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_538_en & cosLUT_MPORT_538_mask) begin
      cosLUT[cosLUT_MPORT_538_addr] <= cosLUT_MPORT_538_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_539_en & cosLUT_MPORT_539_mask) begin
      cosLUT[cosLUT_MPORT_539_addr] <= cosLUT_MPORT_539_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_540_en & cosLUT_MPORT_540_mask) begin
      cosLUT[cosLUT_MPORT_540_addr] <= cosLUT_MPORT_540_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_541_en & cosLUT_MPORT_541_mask) begin
      cosLUT[cosLUT_MPORT_541_addr] <= cosLUT_MPORT_541_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_542_en & cosLUT_MPORT_542_mask) begin
      cosLUT[cosLUT_MPORT_542_addr] <= cosLUT_MPORT_542_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_543_en & cosLUT_MPORT_543_mask) begin
      cosLUT[cosLUT_MPORT_543_addr] <= cosLUT_MPORT_543_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_544_en & cosLUT_MPORT_544_mask) begin
      cosLUT[cosLUT_MPORT_544_addr] <= cosLUT_MPORT_544_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_545_en & cosLUT_MPORT_545_mask) begin
      cosLUT[cosLUT_MPORT_545_addr] <= cosLUT_MPORT_545_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_546_en & cosLUT_MPORT_546_mask) begin
      cosLUT[cosLUT_MPORT_546_addr] <= cosLUT_MPORT_546_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_547_en & cosLUT_MPORT_547_mask) begin
      cosLUT[cosLUT_MPORT_547_addr] <= cosLUT_MPORT_547_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_548_en & cosLUT_MPORT_548_mask) begin
      cosLUT[cosLUT_MPORT_548_addr] <= cosLUT_MPORT_548_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_549_en & cosLUT_MPORT_549_mask) begin
      cosLUT[cosLUT_MPORT_549_addr] <= cosLUT_MPORT_549_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_550_en & cosLUT_MPORT_550_mask) begin
      cosLUT[cosLUT_MPORT_550_addr] <= cosLUT_MPORT_550_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_551_en & cosLUT_MPORT_551_mask) begin
      cosLUT[cosLUT_MPORT_551_addr] <= cosLUT_MPORT_551_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_552_en & cosLUT_MPORT_552_mask) begin
      cosLUT[cosLUT_MPORT_552_addr] <= cosLUT_MPORT_552_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_553_en & cosLUT_MPORT_553_mask) begin
      cosLUT[cosLUT_MPORT_553_addr] <= cosLUT_MPORT_553_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_554_en & cosLUT_MPORT_554_mask) begin
      cosLUT[cosLUT_MPORT_554_addr] <= cosLUT_MPORT_554_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_555_en & cosLUT_MPORT_555_mask) begin
      cosLUT[cosLUT_MPORT_555_addr] <= cosLUT_MPORT_555_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_556_en & cosLUT_MPORT_556_mask) begin
      cosLUT[cosLUT_MPORT_556_addr] <= cosLUT_MPORT_556_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_557_en & cosLUT_MPORT_557_mask) begin
      cosLUT[cosLUT_MPORT_557_addr] <= cosLUT_MPORT_557_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_558_en & cosLUT_MPORT_558_mask) begin
      cosLUT[cosLUT_MPORT_558_addr] <= cosLUT_MPORT_558_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_559_en & cosLUT_MPORT_559_mask) begin
      cosLUT[cosLUT_MPORT_559_addr] <= cosLUT_MPORT_559_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_560_en & cosLUT_MPORT_560_mask) begin
      cosLUT[cosLUT_MPORT_560_addr] <= cosLUT_MPORT_560_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_561_en & cosLUT_MPORT_561_mask) begin
      cosLUT[cosLUT_MPORT_561_addr] <= cosLUT_MPORT_561_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_562_en & cosLUT_MPORT_562_mask) begin
      cosLUT[cosLUT_MPORT_562_addr] <= cosLUT_MPORT_562_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_563_en & cosLUT_MPORT_563_mask) begin
      cosLUT[cosLUT_MPORT_563_addr] <= cosLUT_MPORT_563_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_564_en & cosLUT_MPORT_564_mask) begin
      cosLUT[cosLUT_MPORT_564_addr] <= cosLUT_MPORT_564_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_565_en & cosLUT_MPORT_565_mask) begin
      cosLUT[cosLUT_MPORT_565_addr] <= cosLUT_MPORT_565_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_566_en & cosLUT_MPORT_566_mask) begin
      cosLUT[cosLUT_MPORT_566_addr] <= cosLUT_MPORT_566_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_567_en & cosLUT_MPORT_567_mask) begin
      cosLUT[cosLUT_MPORT_567_addr] <= cosLUT_MPORT_567_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_568_en & cosLUT_MPORT_568_mask) begin
      cosLUT[cosLUT_MPORT_568_addr] <= cosLUT_MPORT_568_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_569_en & cosLUT_MPORT_569_mask) begin
      cosLUT[cosLUT_MPORT_569_addr] <= cosLUT_MPORT_569_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_570_en & cosLUT_MPORT_570_mask) begin
      cosLUT[cosLUT_MPORT_570_addr] <= cosLUT_MPORT_570_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_571_en & cosLUT_MPORT_571_mask) begin
      cosLUT[cosLUT_MPORT_571_addr] <= cosLUT_MPORT_571_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_572_en & cosLUT_MPORT_572_mask) begin
      cosLUT[cosLUT_MPORT_572_addr] <= cosLUT_MPORT_572_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_573_en & cosLUT_MPORT_573_mask) begin
      cosLUT[cosLUT_MPORT_573_addr] <= cosLUT_MPORT_573_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_574_en & cosLUT_MPORT_574_mask) begin
      cosLUT[cosLUT_MPORT_574_addr] <= cosLUT_MPORT_574_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_575_en & cosLUT_MPORT_575_mask) begin
      cosLUT[cosLUT_MPORT_575_addr] <= cosLUT_MPORT_575_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_576_en & cosLUT_MPORT_576_mask) begin
      cosLUT[cosLUT_MPORT_576_addr] <= cosLUT_MPORT_576_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_577_en & cosLUT_MPORT_577_mask) begin
      cosLUT[cosLUT_MPORT_577_addr] <= cosLUT_MPORT_577_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_578_en & cosLUT_MPORT_578_mask) begin
      cosLUT[cosLUT_MPORT_578_addr] <= cosLUT_MPORT_578_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_579_en & cosLUT_MPORT_579_mask) begin
      cosLUT[cosLUT_MPORT_579_addr] <= cosLUT_MPORT_579_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_580_en & cosLUT_MPORT_580_mask) begin
      cosLUT[cosLUT_MPORT_580_addr] <= cosLUT_MPORT_580_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_581_en & cosLUT_MPORT_581_mask) begin
      cosLUT[cosLUT_MPORT_581_addr] <= cosLUT_MPORT_581_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_582_en & cosLUT_MPORT_582_mask) begin
      cosLUT[cosLUT_MPORT_582_addr] <= cosLUT_MPORT_582_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_583_en & cosLUT_MPORT_583_mask) begin
      cosLUT[cosLUT_MPORT_583_addr] <= cosLUT_MPORT_583_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_584_en & cosLUT_MPORT_584_mask) begin
      cosLUT[cosLUT_MPORT_584_addr] <= cosLUT_MPORT_584_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_585_en & cosLUT_MPORT_585_mask) begin
      cosLUT[cosLUT_MPORT_585_addr] <= cosLUT_MPORT_585_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_586_en & cosLUT_MPORT_586_mask) begin
      cosLUT[cosLUT_MPORT_586_addr] <= cosLUT_MPORT_586_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_587_en & cosLUT_MPORT_587_mask) begin
      cosLUT[cosLUT_MPORT_587_addr] <= cosLUT_MPORT_587_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_588_en & cosLUT_MPORT_588_mask) begin
      cosLUT[cosLUT_MPORT_588_addr] <= cosLUT_MPORT_588_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_589_en & cosLUT_MPORT_589_mask) begin
      cosLUT[cosLUT_MPORT_589_addr] <= cosLUT_MPORT_589_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_590_en & cosLUT_MPORT_590_mask) begin
      cosLUT[cosLUT_MPORT_590_addr] <= cosLUT_MPORT_590_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_591_en & cosLUT_MPORT_591_mask) begin
      cosLUT[cosLUT_MPORT_591_addr] <= cosLUT_MPORT_591_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_592_en & cosLUT_MPORT_592_mask) begin
      cosLUT[cosLUT_MPORT_592_addr] <= cosLUT_MPORT_592_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_593_en & cosLUT_MPORT_593_mask) begin
      cosLUT[cosLUT_MPORT_593_addr] <= cosLUT_MPORT_593_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_594_en & cosLUT_MPORT_594_mask) begin
      cosLUT[cosLUT_MPORT_594_addr] <= cosLUT_MPORT_594_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_595_en & cosLUT_MPORT_595_mask) begin
      cosLUT[cosLUT_MPORT_595_addr] <= cosLUT_MPORT_595_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_596_en & cosLUT_MPORT_596_mask) begin
      cosLUT[cosLUT_MPORT_596_addr] <= cosLUT_MPORT_596_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_597_en & cosLUT_MPORT_597_mask) begin
      cosLUT[cosLUT_MPORT_597_addr] <= cosLUT_MPORT_597_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_598_en & cosLUT_MPORT_598_mask) begin
      cosLUT[cosLUT_MPORT_598_addr] <= cosLUT_MPORT_598_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_599_en & cosLUT_MPORT_599_mask) begin
      cosLUT[cosLUT_MPORT_599_addr] <= cosLUT_MPORT_599_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_600_en & cosLUT_MPORT_600_mask) begin
      cosLUT[cosLUT_MPORT_600_addr] <= cosLUT_MPORT_600_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_601_en & cosLUT_MPORT_601_mask) begin
      cosLUT[cosLUT_MPORT_601_addr] <= cosLUT_MPORT_601_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_602_en & cosLUT_MPORT_602_mask) begin
      cosLUT[cosLUT_MPORT_602_addr] <= cosLUT_MPORT_602_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_603_en & cosLUT_MPORT_603_mask) begin
      cosLUT[cosLUT_MPORT_603_addr] <= cosLUT_MPORT_603_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_604_en & cosLUT_MPORT_604_mask) begin
      cosLUT[cosLUT_MPORT_604_addr] <= cosLUT_MPORT_604_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_605_en & cosLUT_MPORT_605_mask) begin
      cosLUT[cosLUT_MPORT_605_addr] <= cosLUT_MPORT_605_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_606_en & cosLUT_MPORT_606_mask) begin
      cosLUT[cosLUT_MPORT_606_addr] <= cosLUT_MPORT_606_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_607_en & cosLUT_MPORT_607_mask) begin
      cosLUT[cosLUT_MPORT_607_addr] <= cosLUT_MPORT_607_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_608_en & cosLUT_MPORT_608_mask) begin
      cosLUT[cosLUT_MPORT_608_addr] <= cosLUT_MPORT_608_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_609_en & cosLUT_MPORT_609_mask) begin
      cosLUT[cosLUT_MPORT_609_addr] <= cosLUT_MPORT_609_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_610_en & cosLUT_MPORT_610_mask) begin
      cosLUT[cosLUT_MPORT_610_addr] <= cosLUT_MPORT_610_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_611_en & cosLUT_MPORT_611_mask) begin
      cosLUT[cosLUT_MPORT_611_addr] <= cosLUT_MPORT_611_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_612_en & cosLUT_MPORT_612_mask) begin
      cosLUT[cosLUT_MPORT_612_addr] <= cosLUT_MPORT_612_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_613_en & cosLUT_MPORT_613_mask) begin
      cosLUT[cosLUT_MPORT_613_addr] <= cosLUT_MPORT_613_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_614_en & cosLUT_MPORT_614_mask) begin
      cosLUT[cosLUT_MPORT_614_addr] <= cosLUT_MPORT_614_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_615_en & cosLUT_MPORT_615_mask) begin
      cosLUT[cosLUT_MPORT_615_addr] <= cosLUT_MPORT_615_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_616_en & cosLUT_MPORT_616_mask) begin
      cosLUT[cosLUT_MPORT_616_addr] <= cosLUT_MPORT_616_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_617_en & cosLUT_MPORT_617_mask) begin
      cosLUT[cosLUT_MPORT_617_addr] <= cosLUT_MPORT_617_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_618_en & cosLUT_MPORT_618_mask) begin
      cosLUT[cosLUT_MPORT_618_addr] <= cosLUT_MPORT_618_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_619_en & cosLUT_MPORT_619_mask) begin
      cosLUT[cosLUT_MPORT_619_addr] <= cosLUT_MPORT_619_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_620_en & cosLUT_MPORT_620_mask) begin
      cosLUT[cosLUT_MPORT_620_addr] <= cosLUT_MPORT_620_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_621_en & cosLUT_MPORT_621_mask) begin
      cosLUT[cosLUT_MPORT_621_addr] <= cosLUT_MPORT_621_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_622_en & cosLUT_MPORT_622_mask) begin
      cosLUT[cosLUT_MPORT_622_addr] <= cosLUT_MPORT_622_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_623_en & cosLUT_MPORT_623_mask) begin
      cosLUT[cosLUT_MPORT_623_addr] <= cosLUT_MPORT_623_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_624_en & cosLUT_MPORT_624_mask) begin
      cosLUT[cosLUT_MPORT_624_addr] <= cosLUT_MPORT_624_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_625_en & cosLUT_MPORT_625_mask) begin
      cosLUT[cosLUT_MPORT_625_addr] <= cosLUT_MPORT_625_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_626_en & cosLUT_MPORT_626_mask) begin
      cosLUT[cosLUT_MPORT_626_addr] <= cosLUT_MPORT_626_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_627_en & cosLUT_MPORT_627_mask) begin
      cosLUT[cosLUT_MPORT_627_addr] <= cosLUT_MPORT_627_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_628_en & cosLUT_MPORT_628_mask) begin
      cosLUT[cosLUT_MPORT_628_addr] <= cosLUT_MPORT_628_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_629_en & cosLUT_MPORT_629_mask) begin
      cosLUT[cosLUT_MPORT_629_addr] <= cosLUT_MPORT_629_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_630_en & cosLUT_MPORT_630_mask) begin
      cosLUT[cosLUT_MPORT_630_addr] <= cosLUT_MPORT_630_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_631_en & cosLUT_MPORT_631_mask) begin
      cosLUT[cosLUT_MPORT_631_addr] <= cosLUT_MPORT_631_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_632_en & cosLUT_MPORT_632_mask) begin
      cosLUT[cosLUT_MPORT_632_addr] <= cosLUT_MPORT_632_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_633_en & cosLUT_MPORT_633_mask) begin
      cosLUT[cosLUT_MPORT_633_addr] <= cosLUT_MPORT_633_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_634_en & cosLUT_MPORT_634_mask) begin
      cosLUT[cosLUT_MPORT_634_addr] <= cosLUT_MPORT_634_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_635_en & cosLUT_MPORT_635_mask) begin
      cosLUT[cosLUT_MPORT_635_addr] <= cosLUT_MPORT_635_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_636_en & cosLUT_MPORT_636_mask) begin
      cosLUT[cosLUT_MPORT_636_addr] <= cosLUT_MPORT_636_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_637_en & cosLUT_MPORT_637_mask) begin
      cosLUT[cosLUT_MPORT_637_addr] <= cosLUT_MPORT_637_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_638_en & cosLUT_MPORT_638_mask) begin
      cosLUT[cosLUT_MPORT_638_addr] <= cosLUT_MPORT_638_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_639_en & cosLUT_MPORT_639_mask) begin
      cosLUT[cosLUT_MPORT_639_addr] <= cosLUT_MPORT_639_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_640_en & cosLUT_MPORT_640_mask) begin
      cosLUT[cosLUT_MPORT_640_addr] <= cosLUT_MPORT_640_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_641_en & cosLUT_MPORT_641_mask) begin
      cosLUT[cosLUT_MPORT_641_addr] <= cosLUT_MPORT_641_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_642_en & cosLUT_MPORT_642_mask) begin
      cosLUT[cosLUT_MPORT_642_addr] <= cosLUT_MPORT_642_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_643_en & cosLUT_MPORT_643_mask) begin
      cosLUT[cosLUT_MPORT_643_addr] <= cosLUT_MPORT_643_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_644_en & cosLUT_MPORT_644_mask) begin
      cosLUT[cosLUT_MPORT_644_addr] <= cosLUT_MPORT_644_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_645_en & cosLUT_MPORT_645_mask) begin
      cosLUT[cosLUT_MPORT_645_addr] <= cosLUT_MPORT_645_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_646_en & cosLUT_MPORT_646_mask) begin
      cosLUT[cosLUT_MPORT_646_addr] <= cosLUT_MPORT_646_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_647_en & cosLUT_MPORT_647_mask) begin
      cosLUT[cosLUT_MPORT_647_addr] <= cosLUT_MPORT_647_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_648_en & cosLUT_MPORT_648_mask) begin
      cosLUT[cosLUT_MPORT_648_addr] <= cosLUT_MPORT_648_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_649_en & cosLUT_MPORT_649_mask) begin
      cosLUT[cosLUT_MPORT_649_addr] <= cosLUT_MPORT_649_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_650_en & cosLUT_MPORT_650_mask) begin
      cosLUT[cosLUT_MPORT_650_addr] <= cosLUT_MPORT_650_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_651_en & cosLUT_MPORT_651_mask) begin
      cosLUT[cosLUT_MPORT_651_addr] <= cosLUT_MPORT_651_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_652_en & cosLUT_MPORT_652_mask) begin
      cosLUT[cosLUT_MPORT_652_addr] <= cosLUT_MPORT_652_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_653_en & cosLUT_MPORT_653_mask) begin
      cosLUT[cosLUT_MPORT_653_addr] <= cosLUT_MPORT_653_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_654_en & cosLUT_MPORT_654_mask) begin
      cosLUT[cosLUT_MPORT_654_addr] <= cosLUT_MPORT_654_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_655_en & cosLUT_MPORT_655_mask) begin
      cosLUT[cosLUT_MPORT_655_addr] <= cosLUT_MPORT_655_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_656_en & cosLUT_MPORT_656_mask) begin
      cosLUT[cosLUT_MPORT_656_addr] <= cosLUT_MPORT_656_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_657_en & cosLUT_MPORT_657_mask) begin
      cosLUT[cosLUT_MPORT_657_addr] <= cosLUT_MPORT_657_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_658_en & cosLUT_MPORT_658_mask) begin
      cosLUT[cosLUT_MPORT_658_addr] <= cosLUT_MPORT_658_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_659_en & cosLUT_MPORT_659_mask) begin
      cosLUT[cosLUT_MPORT_659_addr] <= cosLUT_MPORT_659_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_660_en & cosLUT_MPORT_660_mask) begin
      cosLUT[cosLUT_MPORT_660_addr] <= cosLUT_MPORT_660_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_661_en & cosLUT_MPORT_661_mask) begin
      cosLUT[cosLUT_MPORT_661_addr] <= cosLUT_MPORT_661_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_662_en & cosLUT_MPORT_662_mask) begin
      cosLUT[cosLUT_MPORT_662_addr] <= cosLUT_MPORT_662_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_663_en & cosLUT_MPORT_663_mask) begin
      cosLUT[cosLUT_MPORT_663_addr] <= cosLUT_MPORT_663_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_664_en & cosLUT_MPORT_664_mask) begin
      cosLUT[cosLUT_MPORT_664_addr] <= cosLUT_MPORT_664_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_665_en & cosLUT_MPORT_665_mask) begin
      cosLUT[cosLUT_MPORT_665_addr] <= cosLUT_MPORT_665_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_666_en & cosLUT_MPORT_666_mask) begin
      cosLUT[cosLUT_MPORT_666_addr] <= cosLUT_MPORT_666_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_667_en & cosLUT_MPORT_667_mask) begin
      cosLUT[cosLUT_MPORT_667_addr] <= cosLUT_MPORT_667_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_668_en & cosLUT_MPORT_668_mask) begin
      cosLUT[cosLUT_MPORT_668_addr] <= cosLUT_MPORT_668_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_669_en & cosLUT_MPORT_669_mask) begin
      cosLUT[cosLUT_MPORT_669_addr] <= cosLUT_MPORT_669_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_670_en & cosLUT_MPORT_670_mask) begin
      cosLUT[cosLUT_MPORT_670_addr] <= cosLUT_MPORT_670_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_671_en & cosLUT_MPORT_671_mask) begin
      cosLUT[cosLUT_MPORT_671_addr] <= cosLUT_MPORT_671_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_672_en & cosLUT_MPORT_672_mask) begin
      cosLUT[cosLUT_MPORT_672_addr] <= cosLUT_MPORT_672_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_673_en & cosLUT_MPORT_673_mask) begin
      cosLUT[cosLUT_MPORT_673_addr] <= cosLUT_MPORT_673_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_674_en & cosLUT_MPORT_674_mask) begin
      cosLUT[cosLUT_MPORT_674_addr] <= cosLUT_MPORT_674_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_675_en & cosLUT_MPORT_675_mask) begin
      cosLUT[cosLUT_MPORT_675_addr] <= cosLUT_MPORT_675_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_676_en & cosLUT_MPORT_676_mask) begin
      cosLUT[cosLUT_MPORT_676_addr] <= cosLUT_MPORT_676_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_677_en & cosLUT_MPORT_677_mask) begin
      cosLUT[cosLUT_MPORT_677_addr] <= cosLUT_MPORT_677_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_678_en & cosLUT_MPORT_678_mask) begin
      cosLUT[cosLUT_MPORT_678_addr] <= cosLUT_MPORT_678_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_679_en & cosLUT_MPORT_679_mask) begin
      cosLUT[cosLUT_MPORT_679_addr] <= cosLUT_MPORT_679_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_680_en & cosLUT_MPORT_680_mask) begin
      cosLUT[cosLUT_MPORT_680_addr] <= cosLUT_MPORT_680_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_681_en & cosLUT_MPORT_681_mask) begin
      cosLUT[cosLUT_MPORT_681_addr] <= cosLUT_MPORT_681_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_682_en & cosLUT_MPORT_682_mask) begin
      cosLUT[cosLUT_MPORT_682_addr] <= cosLUT_MPORT_682_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_683_en & cosLUT_MPORT_683_mask) begin
      cosLUT[cosLUT_MPORT_683_addr] <= cosLUT_MPORT_683_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_684_en & cosLUT_MPORT_684_mask) begin
      cosLUT[cosLUT_MPORT_684_addr] <= cosLUT_MPORT_684_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_685_en & cosLUT_MPORT_685_mask) begin
      cosLUT[cosLUT_MPORT_685_addr] <= cosLUT_MPORT_685_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_686_en & cosLUT_MPORT_686_mask) begin
      cosLUT[cosLUT_MPORT_686_addr] <= cosLUT_MPORT_686_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_687_en & cosLUT_MPORT_687_mask) begin
      cosLUT[cosLUT_MPORT_687_addr] <= cosLUT_MPORT_687_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_688_en & cosLUT_MPORT_688_mask) begin
      cosLUT[cosLUT_MPORT_688_addr] <= cosLUT_MPORT_688_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_689_en & cosLUT_MPORT_689_mask) begin
      cosLUT[cosLUT_MPORT_689_addr] <= cosLUT_MPORT_689_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_690_en & cosLUT_MPORT_690_mask) begin
      cosLUT[cosLUT_MPORT_690_addr] <= cosLUT_MPORT_690_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_691_en & cosLUT_MPORT_691_mask) begin
      cosLUT[cosLUT_MPORT_691_addr] <= cosLUT_MPORT_691_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_692_en & cosLUT_MPORT_692_mask) begin
      cosLUT[cosLUT_MPORT_692_addr] <= cosLUT_MPORT_692_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_693_en & cosLUT_MPORT_693_mask) begin
      cosLUT[cosLUT_MPORT_693_addr] <= cosLUT_MPORT_693_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_694_en & cosLUT_MPORT_694_mask) begin
      cosLUT[cosLUT_MPORT_694_addr] <= cosLUT_MPORT_694_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_695_en & cosLUT_MPORT_695_mask) begin
      cosLUT[cosLUT_MPORT_695_addr] <= cosLUT_MPORT_695_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_696_en & cosLUT_MPORT_696_mask) begin
      cosLUT[cosLUT_MPORT_696_addr] <= cosLUT_MPORT_696_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_697_en & cosLUT_MPORT_697_mask) begin
      cosLUT[cosLUT_MPORT_697_addr] <= cosLUT_MPORT_697_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_698_en & cosLUT_MPORT_698_mask) begin
      cosLUT[cosLUT_MPORT_698_addr] <= cosLUT_MPORT_698_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_699_en & cosLUT_MPORT_699_mask) begin
      cosLUT[cosLUT_MPORT_699_addr] <= cosLUT_MPORT_699_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_700_en & cosLUT_MPORT_700_mask) begin
      cosLUT[cosLUT_MPORT_700_addr] <= cosLUT_MPORT_700_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_701_en & cosLUT_MPORT_701_mask) begin
      cosLUT[cosLUT_MPORT_701_addr] <= cosLUT_MPORT_701_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_702_en & cosLUT_MPORT_702_mask) begin
      cosLUT[cosLUT_MPORT_702_addr] <= cosLUT_MPORT_702_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_703_en & cosLUT_MPORT_703_mask) begin
      cosLUT[cosLUT_MPORT_703_addr] <= cosLUT_MPORT_703_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_704_en & cosLUT_MPORT_704_mask) begin
      cosLUT[cosLUT_MPORT_704_addr] <= cosLUT_MPORT_704_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_705_en & cosLUT_MPORT_705_mask) begin
      cosLUT[cosLUT_MPORT_705_addr] <= cosLUT_MPORT_705_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_706_en & cosLUT_MPORT_706_mask) begin
      cosLUT[cosLUT_MPORT_706_addr] <= cosLUT_MPORT_706_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_707_en & cosLUT_MPORT_707_mask) begin
      cosLUT[cosLUT_MPORT_707_addr] <= cosLUT_MPORT_707_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_708_en & cosLUT_MPORT_708_mask) begin
      cosLUT[cosLUT_MPORT_708_addr] <= cosLUT_MPORT_708_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_709_en & cosLUT_MPORT_709_mask) begin
      cosLUT[cosLUT_MPORT_709_addr] <= cosLUT_MPORT_709_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_710_en & cosLUT_MPORT_710_mask) begin
      cosLUT[cosLUT_MPORT_710_addr] <= cosLUT_MPORT_710_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_711_en & cosLUT_MPORT_711_mask) begin
      cosLUT[cosLUT_MPORT_711_addr] <= cosLUT_MPORT_711_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_712_en & cosLUT_MPORT_712_mask) begin
      cosLUT[cosLUT_MPORT_712_addr] <= cosLUT_MPORT_712_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_713_en & cosLUT_MPORT_713_mask) begin
      cosLUT[cosLUT_MPORT_713_addr] <= cosLUT_MPORT_713_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_714_en & cosLUT_MPORT_714_mask) begin
      cosLUT[cosLUT_MPORT_714_addr] <= cosLUT_MPORT_714_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_715_en & cosLUT_MPORT_715_mask) begin
      cosLUT[cosLUT_MPORT_715_addr] <= cosLUT_MPORT_715_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_716_en & cosLUT_MPORT_716_mask) begin
      cosLUT[cosLUT_MPORT_716_addr] <= cosLUT_MPORT_716_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_717_en & cosLUT_MPORT_717_mask) begin
      cosLUT[cosLUT_MPORT_717_addr] <= cosLUT_MPORT_717_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_718_en & cosLUT_MPORT_718_mask) begin
      cosLUT[cosLUT_MPORT_718_addr] <= cosLUT_MPORT_718_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_719_en & cosLUT_MPORT_719_mask) begin
      cosLUT[cosLUT_MPORT_719_addr] <= cosLUT_MPORT_719_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_720_en & cosLUT_MPORT_720_mask) begin
      cosLUT[cosLUT_MPORT_720_addr] <= cosLUT_MPORT_720_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_721_en & cosLUT_MPORT_721_mask) begin
      cosLUT[cosLUT_MPORT_721_addr] <= cosLUT_MPORT_721_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_722_en & cosLUT_MPORT_722_mask) begin
      cosLUT[cosLUT_MPORT_722_addr] <= cosLUT_MPORT_722_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_723_en & cosLUT_MPORT_723_mask) begin
      cosLUT[cosLUT_MPORT_723_addr] <= cosLUT_MPORT_723_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_724_en & cosLUT_MPORT_724_mask) begin
      cosLUT[cosLUT_MPORT_724_addr] <= cosLUT_MPORT_724_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_725_en & cosLUT_MPORT_725_mask) begin
      cosLUT[cosLUT_MPORT_725_addr] <= cosLUT_MPORT_725_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_726_en & cosLUT_MPORT_726_mask) begin
      cosLUT[cosLUT_MPORT_726_addr] <= cosLUT_MPORT_726_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_727_en & cosLUT_MPORT_727_mask) begin
      cosLUT[cosLUT_MPORT_727_addr] <= cosLUT_MPORT_727_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_728_en & cosLUT_MPORT_728_mask) begin
      cosLUT[cosLUT_MPORT_728_addr] <= cosLUT_MPORT_728_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_729_en & cosLUT_MPORT_729_mask) begin
      cosLUT[cosLUT_MPORT_729_addr] <= cosLUT_MPORT_729_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_730_en & cosLUT_MPORT_730_mask) begin
      cosLUT[cosLUT_MPORT_730_addr] <= cosLUT_MPORT_730_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_731_en & cosLUT_MPORT_731_mask) begin
      cosLUT[cosLUT_MPORT_731_addr] <= cosLUT_MPORT_731_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_732_en & cosLUT_MPORT_732_mask) begin
      cosLUT[cosLUT_MPORT_732_addr] <= cosLUT_MPORT_732_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_733_en & cosLUT_MPORT_733_mask) begin
      cosLUT[cosLUT_MPORT_733_addr] <= cosLUT_MPORT_733_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_734_en & cosLUT_MPORT_734_mask) begin
      cosLUT[cosLUT_MPORT_734_addr] <= cosLUT_MPORT_734_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_735_en & cosLUT_MPORT_735_mask) begin
      cosLUT[cosLUT_MPORT_735_addr] <= cosLUT_MPORT_735_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_736_en & cosLUT_MPORT_736_mask) begin
      cosLUT[cosLUT_MPORT_736_addr] <= cosLUT_MPORT_736_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_737_en & cosLUT_MPORT_737_mask) begin
      cosLUT[cosLUT_MPORT_737_addr] <= cosLUT_MPORT_737_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_738_en & cosLUT_MPORT_738_mask) begin
      cosLUT[cosLUT_MPORT_738_addr] <= cosLUT_MPORT_738_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_739_en & cosLUT_MPORT_739_mask) begin
      cosLUT[cosLUT_MPORT_739_addr] <= cosLUT_MPORT_739_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_740_en & cosLUT_MPORT_740_mask) begin
      cosLUT[cosLUT_MPORT_740_addr] <= cosLUT_MPORT_740_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_741_en & cosLUT_MPORT_741_mask) begin
      cosLUT[cosLUT_MPORT_741_addr] <= cosLUT_MPORT_741_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_742_en & cosLUT_MPORT_742_mask) begin
      cosLUT[cosLUT_MPORT_742_addr] <= cosLUT_MPORT_742_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_743_en & cosLUT_MPORT_743_mask) begin
      cosLUT[cosLUT_MPORT_743_addr] <= cosLUT_MPORT_743_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_744_en & cosLUT_MPORT_744_mask) begin
      cosLUT[cosLUT_MPORT_744_addr] <= cosLUT_MPORT_744_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_745_en & cosLUT_MPORT_745_mask) begin
      cosLUT[cosLUT_MPORT_745_addr] <= cosLUT_MPORT_745_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_746_en & cosLUT_MPORT_746_mask) begin
      cosLUT[cosLUT_MPORT_746_addr] <= cosLUT_MPORT_746_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_747_en & cosLUT_MPORT_747_mask) begin
      cosLUT[cosLUT_MPORT_747_addr] <= cosLUT_MPORT_747_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_748_en & cosLUT_MPORT_748_mask) begin
      cosLUT[cosLUT_MPORT_748_addr] <= cosLUT_MPORT_748_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_749_en & cosLUT_MPORT_749_mask) begin
      cosLUT[cosLUT_MPORT_749_addr] <= cosLUT_MPORT_749_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_750_en & cosLUT_MPORT_750_mask) begin
      cosLUT[cosLUT_MPORT_750_addr] <= cosLUT_MPORT_750_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_751_en & cosLUT_MPORT_751_mask) begin
      cosLUT[cosLUT_MPORT_751_addr] <= cosLUT_MPORT_751_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_752_en & cosLUT_MPORT_752_mask) begin
      cosLUT[cosLUT_MPORT_752_addr] <= cosLUT_MPORT_752_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_753_en & cosLUT_MPORT_753_mask) begin
      cosLUT[cosLUT_MPORT_753_addr] <= cosLUT_MPORT_753_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_754_en & cosLUT_MPORT_754_mask) begin
      cosLUT[cosLUT_MPORT_754_addr] <= cosLUT_MPORT_754_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_755_en & cosLUT_MPORT_755_mask) begin
      cosLUT[cosLUT_MPORT_755_addr] <= cosLUT_MPORT_755_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_756_en & cosLUT_MPORT_756_mask) begin
      cosLUT[cosLUT_MPORT_756_addr] <= cosLUT_MPORT_756_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_757_en & cosLUT_MPORT_757_mask) begin
      cosLUT[cosLUT_MPORT_757_addr] <= cosLUT_MPORT_757_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_758_en & cosLUT_MPORT_758_mask) begin
      cosLUT[cosLUT_MPORT_758_addr] <= cosLUT_MPORT_758_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_759_en & cosLUT_MPORT_759_mask) begin
      cosLUT[cosLUT_MPORT_759_addr] <= cosLUT_MPORT_759_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_760_en & cosLUT_MPORT_760_mask) begin
      cosLUT[cosLUT_MPORT_760_addr] <= cosLUT_MPORT_760_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_761_en & cosLUT_MPORT_761_mask) begin
      cosLUT[cosLUT_MPORT_761_addr] <= cosLUT_MPORT_761_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_762_en & cosLUT_MPORT_762_mask) begin
      cosLUT[cosLUT_MPORT_762_addr] <= cosLUT_MPORT_762_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_763_en & cosLUT_MPORT_763_mask) begin
      cosLUT[cosLUT_MPORT_763_addr] <= cosLUT_MPORT_763_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_764_en & cosLUT_MPORT_764_mask) begin
      cosLUT[cosLUT_MPORT_764_addr] <= cosLUT_MPORT_764_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_765_en & cosLUT_MPORT_765_mask) begin
      cosLUT[cosLUT_MPORT_765_addr] <= cosLUT_MPORT_765_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_766_en & cosLUT_MPORT_766_mask) begin
      cosLUT[cosLUT_MPORT_766_addr] <= cosLUT_MPORT_766_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_767_en & cosLUT_MPORT_767_mask) begin
      cosLUT[cosLUT_MPORT_767_addr] <= cosLUT_MPORT_767_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_768_en & cosLUT_MPORT_768_mask) begin
      cosLUT[cosLUT_MPORT_768_addr] <= cosLUT_MPORT_768_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_769_en & cosLUT_MPORT_769_mask) begin
      cosLUT[cosLUT_MPORT_769_addr] <= cosLUT_MPORT_769_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_770_en & cosLUT_MPORT_770_mask) begin
      cosLUT[cosLUT_MPORT_770_addr] <= cosLUT_MPORT_770_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_771_en & cosLUT_MPORT_771_mask) begin
      cosLUT[cosLUT_MPORT_771_addr] <= cosLUT_MPORT_771_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_772_en & cosLUT_MPORT_772_mask) begin
      cosLUT[cosLUT_MPORT_772_addr] <= cosLUT_MPORT_772_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_773_en & cosLUT_MPORT_773_mask) begin
      cosLUT[cosLUT_MPORT_773_addr] <= cosLUT_MPORT_773_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_774_en & cosLUT_MPORT_774_mask) begin
      cosLUT[cosLUT_MPORT_774_addr] <= cosLUT_MPORT_774_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_775_en & cosLUT_MPORT_775_mask) begin
      cosLUT[cosLUT_MPORT_775_addr] <= cosLUT_MPORT_775_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_776_en & cosLUT_MPORT_776_mask) begin
      cosLUT[cosLUT_MPORT_776_addr] <= cosLUT_MPORT_776_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_777_en & cosLUT_MPORT_777_mask) begin
      cosLUT[cosLUT_MPORT_777_addr] <= cosLUT_MPORT_777_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_778_en & cosLUT_MPORT_778_mask) begin
      cosLUT[cosLUT_MPORT_778_addr] <= cosLUT_MPORT_778_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_779_en & cosLUT_MPORT_779_mask) begin
      cosLUT[cosLUT_MPORT_779_addr] <= cosLUT_MPORT_779_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_780_en & cosLUT_MPORT_780_mask) begin
      cosLUT[cosLUT_MPORT_780_addr] <= cosLUT_MPORT_780_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_781_en & cosLUT_MPORT_781_mask) begin
      cosLUT[cosLUT_MPORT_781_addr] <= cosLUT_MPORT_781_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_782_en & cosLUT_MPORT_782_mask) begin
      cosLUT[cosLUT_MPORT_782_addr] <= cosLUT_MPORT_782_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_783_en & cosLUT_MPORT_783_mask) begin
      cosLUT[cosLUT_MPORT_783_addr] <= cosLUT_MPORT_783_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_784_en & cosLUT_MPORT_784_mask) begin
      cosLUT[cosLUT_MPORT_784_addr] <= cosLUT_MPORT_784_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_785_en & cosLUT_MPORT_785_mask) begin
      cosLUT[cosLUT_MPORT_785_addr] <= cosLUT_MPORT_785_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_786_en & cosLUT_MPORT_786_mask) begin
      cosLUT[cosLUT_MPORT_786_addr] <= cosLUT_MPORT_786_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_787_en & cosLUT_MPORT_787_mask) begin
      cosLUT[cosLUT_MPORT_787_addr] <= cosLUT_MPORT_787_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_788_en & cosLUT_MPORT_788_mask) begin
      cosLUT[cosLUT_MPORT_788_addr] <= cosLUT_MPORT_788_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_789_en & cosLUT_MPORT_789_mask) begin
      cosLUT[cosLUT_MPORT_789_addr] <= cosLUT_MPORT_789_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_790_en & cosLUT_MPORT_790_mask) begin
      cosLUT[cosLUT_MPORT_790_addr] <= cosLUT_MPORT_790_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_791_en & cosLUT_MPORT_791_mask) begin
      cosLUT[cosLUT_MPORT_791_addr] <= cosLUT_MPORT_791_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_792_en & cosLUT_MPORT_792_mask) begin
      cosLUT[cosLUT_MPORT_792_addr] <= cosLUT_MPORT_792_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_793_en & cosLUT_MPORT_793_mask) begin
      cosLUT[cosLUT_MPORT_793_addr] <= cosLUT_MPORT_793_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_794_en & cosLUT_MPORT_794_mask) begin
      cosLUT[cosLUT_MPORT_794_addr] <= cosLUT_MPORT_794_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_795_en & cosLUT_MPORT_795_mask) begin
      cosLUT[cosLUT_MPORT_795_addr] <= cosLUT_MPORT_795_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_796_en & cosLUT_MPORT_796_mask) begin
      cosLUT[cosLUT_MPORT_796_addr] <= cosLUT_MPORT_796_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_797_en & cosLUT_MPORT_797_mask) begin
      cosLUT[cosLUT_MPORT_797_addr] <= cosLUT_MPORT_797_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_798_en & cosLUT_MPORT_798_mask) begin
      cosLUT[cosLUT_MPORT_798_addr] <= cosLUT_MPORT_798_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_799_en & cosLUT_MPORT_799_mask) begin
      cosLUT[cosLUT_MPORT_799_addr] <= cosLUT_MPORT_799_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_800_en & cosLUT_MPORT_800_mask) begin
      cosLUT[cosLUT_MPORT_800_addr] <= cosLUT_MPORT_800_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_801_en & cosLUT_MPORT_801_mask) begin
      cosLUT[cosLUT_MPORT_801_addr] <= cosLUT_MPORT_801_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_802_en & cosLUT_MPORT_802_mask) begin
      cosLUT[cosLUT_MPORT_802_addr] <= cosLUT_MPORT_802_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_803_en & cosLUT_MPORT_803_mask) begin
      cosLUT[cosLUT_MPORT_803_addr] <= cosLUT_MPORT_803_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_804_en & cosLUT_MPORT_804_mask) begin
      cosLUT[cosLUT_MPORT_804_addr] <= cosLUT_MPORT_804_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_805_en & cosLUT_MPORT_805_mask) begin
      cosLUT[cosLUT_MPORT_805_addr] <= cosLUT_MPORT_805_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_806_en & cosLUT_MPORT_806_mask) begin
      cosLUT[cosLUT_MPORT_806_addr] <= cosLUT_MPORT_806_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_807_en & cosLUT_MPORT_807_mask) begin
      cosLUT[cosLUT_MPORT_807_addr] <= cosLUT_MPORT_807_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_808_en & cosLUT_MPORT_808_mask) begin
      cosLUT[cosLUT_MPORT_808_addr] <= cosLUT_MPORT_808_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_809_en & cosLUT_MPORT_809_mask) begin
      cosLUT[cosLUT_MPORT_809_addr] <= cosLUT_MPORT_809_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_810_en & cosLUT_MPORT_810_mask) begin
      cosLUT[cosLUT_MPORT_810_addr] <= cosLUT_MPORT_810_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_811_en & cosLUT_MPORT_811_mask) begin
      cosLUT[cosLUT_MPORT_811_addr] <= cosLUT_MPORT_811_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_812_en & cosLUT_MPORT_812_mask) begin
      cosLUT[cosLUT_MPORT_812_addr] <= cosLUT_MPORT_812_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_813_en & cosLUT_MPORT_813_mask) begin
      cosLUT[cosLUT_MPORT_813_addr] <= cosLUT_MPORT_813_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_814_en & cosLUT_MPORT_814_mask) begin
      cosLUT[cosLUT_MPORT_814_addr] <= cosLUT_MPORT_814_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_815_en & cosLUT_MPORT_815_mask) begin
      cosLUT[cosLUT_MPORT_815_addr] <= cosLUT_MPORT_815_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_816_en & cosLUT_MPORT_816_mask) begin
      cosLUT[cosLUT_MPORT_816_addr] <= cosLUT_MPORT_816_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_817_en & cosLUT_MPORT_817_mask) begin
      cosLUT[cosLUT_MPORT_817_addr] <= cosLUT_MPORT_817_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_818_en & cosLUT_MPORT_818_mask) begin
      cosLUT[cosLUT_MPORT_818_addr] <= cosLUT_MPORT_818_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_819_en & cosLUT_MPORT_819_mask) begin
      cosLUT[cosLUT_MPORT_819_addr] <= cosLUT_MPORT_819_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_820_en & cosLUT_MPORT_820_mask) begin
      cosLUT[cosLUT_MPORT_820_addr] <= cosLUT_MPORT_820_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_821_en & cosLUT_MPORT_821_mask) begin
      cosLUT[cosLUT_MPORT_821_addr] <= cosLUT_MPORT_821_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_822_en & cosLUT_MPORT_822_mask) begin
      cosLUT[cosLUT_MPORT_822_addr] <= cosLUT_MPORT_822_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_823_en & cosLUT_MPORT_823_mask) begin
      cosLUT[cosLUT_MPORT_823_addr] <= cosLUT_MPORT_823_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_824_en & cosLUT_MPORT_824_mask) begin
      cosLUT[cosLUT_MPORT_824_addr] <= cosLUT_MPORT_824_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_825_en & cosLUT_MPORT_825_mask) begin
      cosLUT[cosLUT_MPORT_825_addr] <= cosLUT_MPORT_825_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_826_en & cosLUT_MPORT_826_mask) begin
      cosLUT[cosLUT_MPORT_826_addr] <= cosLUT_MPORT_826_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_827_en & cosLUT_MPORT_827_mask) begin
      cosLUT[cosLUT_MPORT_827_addr] <= cosLUT_MPORT_827_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_828_en & cosLUT_MPORT_828_mask) begin
      cosLUT[cosLUT_MPORT_828_addr] <= cosLUT_MPORT_828_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_829_en & cosLUT_MPORT_829_mask) begin
      cosLUT[cosLUT_MPORT_829_addr] <= cosLUT_MPORT_829_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_830_en & cosLUT_MPORT_830_mask) begin
      cosLUT[cosLUT_MPORT_830_addr] <= cosLUT_MPORT_830_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_831_en & cosLUT_MPORT_831_mask) begin
      cosLUT[cosLUT_MPORT_831_addr] <= cosLUT_MPORT_831_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_832_en & cosLUT_MPORT_832_mask) begin
      cosLUT[cosLUT_MPORT_832_addr] <= cosLUT_MPORT_832_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_833_en & cosLUT_MPORT_833_mask) begin
      cosLUT[cosLUT_MPORT_833_addr] <= cosLUT_MPORT_833_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_834_en & cosLUT_MPORT_834_mask) begin
      cosLUT[cosLUT_MPORT_834_addr] <= cosLUT_MPORT_834_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_835_en & cosLUT_MPORT_835_mask) begin
      cosLUT[cosLUT_MPORT_835_addr] <= cosLUT_MPORT_835_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_836_en & cosLUT_MPORT_836_mask) begin
      cosLUT[cosLUT_MPORT_836_addr] <= cosLUT_MPORT_836_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_837_en & cosLUT_MPORT_837_mask) begin
      cosLUT[cosLUT_MPORT_837_addr] <= cosLUT_MPORT_837_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_838_en & cosLUT_MPORT_838_mask) begin
      cosLUT[cosLUT_MPORT_838_addr] <= cosLUT_MPORT_838_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_839_en & cosLUT_MPORT_839_mask) begin
      cosLUT[cosLUT_MPORT_839_addr] <= cosLUT_MPORT_839_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_840_en & cosLUT_MPORT_840_mask) begin
      cosLUT[cosLUT_MPORT_840_addr] <= cosLUT_MPORT_840_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_841_en & cosLUT_MPORT_841_mask) begin
      cosLUT[cosLUT_MPORT_841_addr] <= cosLUT_MPORT_841_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_842_en & cosLUT_MPORT_842_mask) begin
      cosLUT[cosLUT_MPORT_842_addr] <= cosLUT_MPORT_842_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_843_en & cosLUT_MPORT_843_mask) begin
      cosLUT[cosLUT_MPORT_843_addr] <= cosLUT_MPORT_843_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_844_en & cosLUT_MPORT_844_mask) begin
      cosLUT[cosLUT_MPORT_844_addr] <= cosLUT_MPORT_844_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_845_en & cosLUT_MPORT_845_mask) begin
      cosLUT[cosLUT_MPORT_845_addr] <= cosLUT_MPORT_845_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_846_en & cosLUT_MPORT_846_mask) begin
      cosLUT[cosLUT_MPORT_846_addr] <= cosLUT_MPORT_846_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_847_en & cosLUT_MPORT_847_mask) begin
      cosLUT[cosLUT_MPORT_847_addr] <= cosLUT_MPORT_847_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_848_en & cosLUT_MPORT_848_mask) begin
      cosLUT[cosLUT_MPORT_848_addr] <= cosLUT_MPORT_848_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_849_en & cosLUT_MPORT_849_mask) begin
      cosLUT[cosLUT_MPORT_849_addr] <= cosLUT_MPORT_849_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_850_en & cosLUT_MPORT_850_mask) begin
      cosLUT[cosLUT_MPORT_850_addr] <= cosLUT_MPORT_850_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_851_en & cosLUT_MPORT_851_mask) begin
      cosLUT[cosLUT_MPORT_851_addr] <= cosLUT_MPORT_851_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_852_en & cosLUT_MPORT_852_mask) begin
      cosLUT[cosLUT_MPORT_852_addr] <= cosLUT_MPORT_852_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_853_en & cosLUT_MPORT_853_mask) begin
      cosLUT[cosLUT_MPORT_853_addr] <= cosLUT_MPORT_853_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_854_en & cosLUT_MPORT_854_mask) begin
      cosLUT[cosLUT_MPORT_854_addr] <= cosLUT_MPORT_854_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_855_en & cosLUT_MPORT_855_mask) begin
      cosLUT[cosLUT_MPORT_855_addr] <= cosLUT_MPORT_855_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_856_en & cosLUT_MPORT_856_mask) begin
      cosLUT[cosLUT_MPORT_856_addr] <= cosLUT_MPORT_856_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_857_en & cosLUT_MPORT_857_mask) begin
      cosLUT[cosLUT_MPORT_857_addr] <= cosLUT_MPORT_857_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_858_en & cosLUT_MPORT_858_mask) begin
      cosLUT[cosLUT_MPORT_858_addr] <= cosLUT_MPORT_858_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_859_en & cosLUT_MPORT_859_mask) begin
      cosLUT[cosLUT_MPORT_859_addr] <= cosLUT_MPORT_859_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_860_en & cosLUT_MPORT_860_mask) begin
      cosLUT[cosLUT_MPORT_860_addr] <= cosLUT_MPORT_860_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_861_en & cosLUT_MPORT_861_mask) begin
      cosLUT[cosLUT_MPORT_861_addr] <= cosLUT_MPORT_861_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_862_en & cosLUT_MPORT_862_mask) begin
      cosLUT[cosLUT_MPORT_862_addr] <= cosLUT_MPORT_862_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_863_en & cosLUT_MPORT_863_mask) begin
      cosLUT[cosLUT_MPORT_863_addr] <= cosLUT_MPORT_863_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_864_en & cosLUT_MPORT_864_mask) begin
      cosLUT[cosLUT_MPORT_864_addr] <= cosLUT_MPORT_864_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_865_en & cosLUT_MPORT_865_mask) begin
      cosLUT[cosLUT_MPORT_865_addr] <= cosLUT_MPORT_865_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_866_en & cosLUT_MPORT_866_mask) begin
      cosLUT[cosLUT_MPORT_866_addr] <= cosLUT_MPORT_866_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_867_en & cosLUT_MPORT_867_mask) begin
      cosLUT[cosLUT_MPORT_867_addr] <= cosLUT_MPORT_867_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_868_en & cosLUT_MPORT_868_mask) begin
      cosLUT[cosLUT_MPORT_868_addr] <= cosLUT_MPORT_868_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_869_en & cosLUT_MPORT_869_mask) begin
      cosLUT[cosLUT_MPORT_869_addr] <= cosLUT_MPORT_869_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_870_en & cosLUT_MPORT_870_mask) begin
      cosLUT[cosLUT_MPORT_870_addr] <= cosLUT_MPORT_870_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_871_en & cosLUT_MPORT_871_mask) begin
      cosLUT[cosLUT_MPORT_871_addr] <= cosLUT_MPORT_871_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_872_en & cosLUT_MPORT_872_mask) begin
      cosLUT[cosLUT_MPORT_872_addr] <= cosLUT_MPORT_872_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_873_en & cosLUT_MPORT_873_mask) begin
      cosLUT[cosLUT_MPORT_873_addr] <= cosLUT_MPORT_873_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_874_en & cosLUT_MPORT_874_mask) begin
      cosLUT[cosLUT_MPORT_874_addr] <= cosLUT_MPORT_874_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_875_en & cosLUT_MPORT_875_mask) begin
      cosLUT[cosLUT_MPORT_875_addr] <= cosLUT_MPORT_875_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_876_en & cosLUT_MPORT_876_mask) begin
      cosLUT[cosLUT_MPORT_876_addr] <= cosLUT_MPORT_876_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_877_en & cosLUT_MPORT_877_mask) begin
      cosLUT[cosLUT_MPORT_877_addr] <= cosLUT_MPORT_877_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_878_en & cosLUT_MPORT_878_mask) begin
      cosLUT[cosLUT_MPORT_878_addr] <= cosLUT_MPORT_878_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_879_en & cosLUT_MPORT_879_mask) begin
      cosLUT[cosLUT_MPORT_879_addr] <= cosLUT_MPORT_879_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_880_en & cosLUT_MPORT_880_mask) begin
      cosLUT[cosLUT_MPORT_880_addr] <= cosLUT_MPORT_880_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_881_en & cosLUT_MPORT_881_mask) begin
      cosLUT[cosLUT_MPORT_881_addr] <= cosLUT_MPORT_881_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_882_en & cosLUT_MPORT_882_mask) begin
      cosLUT[cosLUT_MPORT_882_addr] <= cosLUT_MPORT_882_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_883_en & cosLUT_MPORT_883_mask) begin
      cosLUT[cosLUT_MPORT_883_addr] <= cosLUT_MPORT_883_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_884_en & cosLUT_MPORT_884_mask) begin
      cosLUT[cosLUT_MPORT_884_addr] <= cosLUT_MPORT_884_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_885_en & cosLUT_MPORT_885_mask) begin
      cosLUT[cosLUT_MPORT_885_addr] <= cosLUT_MPORT_885_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_886_en & cosLUT_MPORT_886_mask) begin
      cosLUT[cosLUT_MPORT_886_addr] <= cosLUT_MPORT_886_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_887_en & cosLUT_MPORT_887_mask) begin
      cosLUT[cosLUT_MPORT_887_addr] <= cosLUT_MPORT_887_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_888_en & cosLUT_MPORT_888_mask) begin
      cosLUT[cosLUT_MPORT_888_addr] <= cosLUT_MPORT_888_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_889_en & cosLUT_MPORT_889_mask) begin
      cosLUT[cosLUT_MPORT_889_addr] <= cosLUT_MPORT_889_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_890_en & cosLUT_MPORT_890_mask) begin
      cosLUT[cosLUT_MPORT_890_addr] <= cosLUT_MPORT_890_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_891_en & cosLUT_MPORT_891_mask) begin
      cosLUT[cosLUT_MPORT_891_addr] <= cosLUT_MPORT_891_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_892_en & cosLUT_MPORT_892_mask) begin
      cosLUT[cosLUT_MPORT_892_addr] <= cosLUT_MPORT_892_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_893_en & cosLUT_MPORT_893_mask) begin
      cosLUT[cosLUT_MPORT_893_addr] <= cosLUT_MPORT_893_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_894_en & cosLUT_MPORT_894_mask) begin
      cosLUT[cosLUT_MPORT_894_addr] <= cosLUT_MPORT_894_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_895_en & cosLUT_MPORT_895_mask) begin
      cosLUT[cosLUT_MPORT_895_addr] <= cosLUT_MPORT_895_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_896_en & cosLUT_MPORT_896_mask) begin
      cosLUT[cosLUT_MPORT_896_addr] <= cosLUT_MPORT_896_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_897_en & cosLUT_MPORT_897_mask) begin
      cosLUT[cosLUT_MPORT_897_addr] <= cosLUT_MPORT_897_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_898_en & cosLUT_MPORT_898_mask) begin
      cosLUT[cosLUT_MPORT_898_addr] <= cosLUT_MPORT_898_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_899_en & cosLUT_MPORT_899_mask) begin
      cosLUT[cosLUT_MPORT_899_addr] <= cosLUT_MPORT_899_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_900_en & cosLUT_MPORT_900_mask) begin
      cosLUT[cosLUT_MPORT_900_addr] <= cosLUT_MPORT_900_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_901_en & cosLUT_MPORT_901_mask) begin
      cosLUT[cosLUT_MPORT_901_addr] <= cosLUT_MPORT_901_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_902_en & cosLUT_MPORT_902_mask) begin
      cosLUT[cosLUT_MPORT_902_addr] <= cosLUT_MPORT_902_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_903_en & cosLUT_MPORT_903_mask) begin
      cosLUT[cosLUT_MPORT_903_addr] <= cosLUT_MPORT_903_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_904_en & cosLUT_MPORT_904_mask) begin
      cosLUT[cosLUT_MPORT_904_addr] <= cosLUT_MPORT_904_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_905_en & cosLUT_MPORT_905_mask) begin
      cosLUT[cosLUT_MPORT_905_addr] <= cosLUT_MPORT_905_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_906_en & cosLUT_MPORT_906_mask) begin
      cosLUT[cosLUT_MPORT_906_addr] <= cosLUT_MPORT_906_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_907_en & cosLUT_MPORT_907_mask) begin
      cosLUT[cosLUT_MPORT_907_addr] <= cosLUT_MPORT_907_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_908_en & cosLUT_MPORT_908_mask) begin
      cosLUT[cosLUT_MPORT_908_addr] <= cosLUT_MPORT_908_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_909_en & cosLUT_MPORT_909_mask) begin
      cosLUT[cosLUT_MPORT_909_addr] <= cosLUT_MPORT_909_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_910_en & cosLUT_MPORT_910_mask) begin
      cosLUT[cosLUT_MPORT_910_addr] <= cosLUT_MPORT_910_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_911_en & cosLUT_MPORT_911_mask) begin
      cosLUT[cosLUT_MPORT_911_addr] <= cosLUT_MPORT_911_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_912_en & cosLUT_MPORT_912_mask) begin
      cosLUT[cosLUT_MPORT_912_addr] <= cosLUT_MPORT_912_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_913_en & cosLUT_MPORT_913_mask) begin
      cosLUT[cosLUT_MPORT_913_addr] <= cosLUT_MPORT_913_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_914_en & cosLUT_MPORT_914_mask) begin
      cosLUT[cosLUT_MPORT_914_addr] <= cosLUT_MPORT_914_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_915_en & cosLUT_MPORT_915_mask) begin
      cosLUT[cosLUT_MPORT_915_addr] <= cosLUT_MPORT_915_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_916_en & cosLUT_MPORT_916_mask) begin
      cosLUT[cosLUT_MPORT_916_addr] <= cosLUT_MPORT_916_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_917_en & cosLUT_MPORT_917_mask) begin
      cosLUT[cosLUT_MPORT_917_addr] <= cosLUT_MPORT_917_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_918_en & cosLUT_MPORT_918_mask) begin
      cosLUT[cosLUT_MPORT_918_addr] <= cosLUT_MPORT_918_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_919_en & cosLUT_MPORT_919_mask) begin
      cosLUT[cosLUT_MPORT_919_addr] <= cosLUT_MPORT_919_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_920_en & cosLUT_MPORT_920_mask) begin
      cosLUT[cosLUT_MPORT_920_addr] <= cosLUT_MPORT_920_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_921_en & cosLUT_MPORT_921_mask) begin
      cosLUT[cosLUT_MPORT_921_addr] <= cosLUT_MPORT_921_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_922_en & cosLUT_MPORT_922_mask) begin
      cosLUT[cosLUT_MPORT_922_addr] <= cosLUT_MPORT_922_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_923_en & cosLUT_MPORT_923_mask) begin
      cosLUT[cosLUT_MPORT_923_addr] <= cosLUT_MPORT_923_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_924_en & cosLUT_MPORT_924_mask) begin
      cosLUT[cosLUT_MPORT_924_addr] <= cosLUT_MPORT_924_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_925_en & cosLUT_MPORT_925_mask) begin
      cosLUT[cosLUT_MPORT_925_addr] <= cosLUT_MPORT_925_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_926_en & cosLUT_MPORT_926_mask) begin
      cosLUT[cosLUT_MPORT_926_addr] <= cosLUT_MPORT_926_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_927_en & cosLUT_MPORT_927_mask) begin
      cosLUT[cosLUT_MPORT_927_addr] <= cosLUT_MPORT_927_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_928_en & cosLUT_MPORT_928_mask) begin
      cosLUT[cosLUT_MPORT_928_addr] <= cosLUT_MPORT_928_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_929_en & cosLUT_MPORT_929_mask) begin
      cosLUT[cosLUT_MPORT_929_addr] <= cosLUT_MPORT_929_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_930_en & cosLUT_MPORT_930_mask) begin
      cosLUT[cosLUT_MPORT_930_addr] <= cosLUT_MPORT_930_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_931_en & cosLUT_MPORT_931_mask) begin
      cosLUT[cosLUT_MPORT_931_addr] <= cosLUT_MPORT_931_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_932_en & cosLUT_MPORT_932_mask) begin
      cosLUT[cosLUT_MPORT_932_addr] <= cosLUT_MPORT_932_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_933_en & cosLUT_MPORT_933_mask) begin
      cosLUT[cosLUT_MPORT_933_addr] <= cosLUT_MPORT_933_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_934_en & cosLUT_MPORT_934_mask) begin
      cosLUT[cosLUT_MPORT_934_addr] <= cosLUT_MPORT_934_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_935_en & cosLUT_MPORT_935_mask) begin
      cosLUT[cosLUT_MPORT_935_addr] <= cosLUT_MPORT_935_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_936_en & cosLUT_MPORT_936_mask) begin
      cosLUT[cosLUT_MPORT_936_addr] <= cosLUT_MPORT_936_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_937_en & cosLUT_MPORT_937_mask) begin
      cosLUT[cosLUT_MPORT_937_addr] <= cosLUT_MPORT_937_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_938_en & cosLUT_MPORT_938_mask) begin
      cosLUT[cosLUT_MPORT_938_addr] <= cosLUT_MPORT_938_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_939_en & cosLUT_MPORT_939_mask) begin
      cosLUT[cosLUT_MPORT_939_addr] <= cosLUT_MPORT_939_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_940_en & cosLUT_MPORT_940_mask) begin
      cosLUT[cosLUT_MPORT_940_addr] <= cosLUT_MPORT_940_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_941_en & cosLUT_MPORT_941_mask) begin
      cosLUT[cosLUT_MPORT_941_addr] <= cosLUT_MPORT_941_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_942_en & cosLUT_MPORT_942_mask) begin
      cosLUT[cosLUT_MPORT_942_addr] <= cosLUT_MPORT_942_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_943_en & cosLUT_MPORT_943_mask) begin
      cosLUT[cosLUT_MPORT_943_addr] <= cosLUT_MPORT_943_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_944_en & cosLUT_MPORT_944_mask) begin
      cosLUT[cosLUT_MPORT_944_addr] <= cosLUT_MPORT_944_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_945_en & cosLUT_MPORT_945_mask) begin
      cosLUT[cosLUT_MPORT_945_addr] <= cosLUT_MPORT_945_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_946_en & cosLUT_MPORT_946_mask) begin
      cosLUT[cosLUT_MPORT_946_addr] <= cosLUT_MPORT_946_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_947_en & cosLUT_MPORT_947_mask) begin
      cosLUT[cosLUT_MPORT_947_addr] <= cosLUT_MPORT_947_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_948_en & cosLUT_MPORT_948_mask) begin
      cosLUT[cosLUT_MPORT_948_addr] <= cosLUT_MPORT_948_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_949_en & cosLUT_MPORT_949_mask) begin
      cosLUT[cosLUT_MPORT_949_addr] <= cosLUT_MPORT_949_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_950_en & cosLUT_MPORT_950_mask) begin
      cosLUT[cosLUT_MPORT_950_addr] <= cosLUT_MPORT_950_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_951_en & cosLUT_MPORT_951_mask) begin
      cosLUT[cosLUT_MPORT_951_addr] <= cosLUT_MPORT_951_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_952_en & cosLUT_MPORT_952_mask) begin
      cosLUT[cosLUT_MPORT_952_addr] <= cosLUT_MPORT_952_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_953_en & cosLUT_MPORT_953_mask) begin
      cosLUT[cosLUT_MPORT_953_addr] <= cosLUT_MPORT_953_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_954_en & cosLUT_MPORT_954_mask) begin
      cosLUT[cosLUT_MPORT_954_addr] <= cosLUT_MPORT_954_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_955_en & cosLUT_MPORT_955_mask) begin
      cosLUT[cosLUT_MPORT_955_addr] <= cosLUT_MPORT_955_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_956_en & cosLUT_MPORT_956_mask) begin
      cosLUT[cosLUT_MPORT_956_addr] <= cosLUT_MPORT_956_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_957_en & cosLUT_MPORT_957_mask) begin
      cosLUT[cosLUT_MPORT_957_addr] <= cosLUT_MPORT_957_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_958_en & cosLUT_MPORT_958_mask) begin
      cosLUT[cosLUT_MPORT_958_addr] <= cosLUT_MPORT_958_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_959_en & cosLUT_MPORT_959_mask) begin
      cosLUT[cosLUT_MPORT_959_addr] <= cosLUT_MPORT_959_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_960_en & cosLUT_MPORT_960_mask) begin
      cosLUT[cosLUT_MPORT_960_addr] <= cosLUT_MPORT_960_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_961_en & cosLUT_MPORT_961_mask) begin
      cosLUT[cosLUT_MPORT_961_addr] <= cosLUT_MPORT_961_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_962_en & cosLUT_MPORT_962_mask) begin
      cosLUT[cosLUT_MPORT_962_addr] <= cosLUT_MPORT_962_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_963_en & cosLUT_MPORT_963_mask) begin
      cosLUT[cosLUT_MPORT_963_addr] <= cosLUT_MPORT_963_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_964_en & cosLUT_MPORT_964_mask) begin
      cosLUT[cosLUT_MPORT_964_addr] <= cosLUT_MPORT_964_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_965_en & cosLUT_MPORT_965_mask) begin
      cosLUT[cosLUT_MPORT_965_addr] <= cosLUT_MPORT_965_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_966_en & cosLUT_MPORT_966_mask) begin
      cosLUT[cosLUT_MPORT_966_addr] <= cosLUT_MPORT_966_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_967_en & cosLUT_MPORT_967_mask) begin
      cosLUT[cosLUT_MPORT_967_addr] <= cosLUT_MPORT_967_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_968_en & cosLUT_MPORT_968_mask) begin
      cosLUT[cosLUT_MPORT_968_addr] <= cosLUT_MPORT_968_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_969_en & cosLUT_MPORT_969_mask) begin
      cosLUT[cosLUT_MPORT_969_addr] <= cosLUT_MPORT_969_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_970_en & cosLUT_MPORT_970_mask) begin
      cosLUT[cosLUT_MPORT_970_addr] <= cosLUT_MPORT_970_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_971_en & cosLUT_MPORT_971_mask) begin
      cosLUT[cosLUT_MPORT_971_addr] <= cosLUT_MPORT_971_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_972_en & cosLUT_MPORT_972_mask) begin
      cosLUT[cosLUT_MPORT_972_addr] <= cosLUT_MPORT_972_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_973_en & cosLUT_MPORT_973_mask) begin
      cosLUT[cosLUT_MPORT_973_addr] <= cosLUT_MPORT_973_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_974_en & cosLUT_MPORT_974_mask) begin
      cosLUT[cosLUT_MPORT_974_addr] <= cosLUT_MPORT_974_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_975_en & cosLUT_MPORT_975_mask) begin
      cosLUT[cosLUT_MPORT_975_addr] <= cosLUT_MPORT_975_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_976_en & cosLUT_MPORT_976_mask) begin
      cosLUT[cosLUT_MPORT_976_addr] <= cosLUT_MPORT_976_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_977_en & cosLUT_MPORT_977_mask) begin
      cosLUT[cosLUT_MPORT_977_addr] <= cosLUT_MPORT_977_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_978_en & cosLUT_MPORT_978_mask) begin
      cosLUT[cosLUT_MPORT_978_addr] <= cosLUT_MPORT_978_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_979_en & cosLUT_MPORT_979_mask) begin
      cosLUT[cosLUT_MPORT_979_addr] <= cosLUT_MPORT_979_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_980_en & cosLUT_MPORT_980_mask) begin
      cosLUT[cosLUT_MPORT_980_addr] <= cosLUT_MPORT_980_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_981_en & cosLUT_MPORT_981_mask) begin
      cosLUT[cosLUT_MPORT_981_addr] <= cosLUT_MPORT_981_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_982_en & cosLUT_MPORT_982_mask) begin
      cosLUT[cosLUT_MPORT_982_addr] <= cosLUT_MPORT_982_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_983_en & cosLUT_MPORT_983_mask) begin
      cosLUT[cosLUT_MPORT_983_addr] <= cosLUT_MPORT_983_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_984_en & cosLUT_MPORT_984_mask) begin
      cosLUT[cosLUT_MPORT_984_addr] <= cosLUT_MPORT_984_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_985_en & cosLUT_MPORT_985_mask) begin
      cosLUT[cosLUT_MPORT_985_addr] <= cosLUT_MPORT_985_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_986_en & cosLUT_MPORT_986_mask) begin
      cosLUT[cosLUT_MPORT_986_addr] <= cosLUT_MPORT_986_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_987_en & cosLUT_MPORT_987_mask) begin
      cosLUT[cosLUT_MPORT_987_addr] <= cosLUT_MPORT_987_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_988_en & cosLUT_MPORT_988_mask) begin
      cosLUT[cosLUT_MPORT_988_addr] <= cosLUT_MPORT_988_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_989_en & cosLUT_MPORT_989_mask) begin
      cosLUT[cosLUT_MPORT_989_addr] <= cosLUT_MPORT_989_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_990_en & cosLUT_MPORT_990_mask) begin
      cosLUT[cosLUT_MPORT_990_addr] <= cosLUT_MPORT_990_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_991_en & cosLUT_MPORT_991_mask) begin
      cosLUT[cosLUT_MPORT_991_addr] <= cosLUT_MPORT_991_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_992_en & cosLUT_MPORT_992_mask) begin
      cosLUT[cosLUT_MPORT_992_addr] <= cosLUT_MPORT_992_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_993_en & cosLUT_MPORT_993_mask) begin
      cosLUT[cosLUT_MPORT_993_addr] <= cosLUT_MPORT_993_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_994_en & cosLUT_MPORT_994_mask) begin
      cosLUT[cosLUT_MPORT_994_addr] <= cosLUT_MPORT_994_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_995_en & cosLUT_MPORT_995_mask) begin
      cosLUT[cosLUT_MPORT_995_addr] <= cosLUT_MPORT_995_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_996_en & cosLUT_MPORT_996_mask) begin
      cosLUT[cosLUT_MPORT_996_addr] <= cosLUT_MPORT_996_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_997_en & cosLUT_MPORT_997_mask) begin
      cosLUT[cosLUT_MPORT_997_addr] <= cosLUT_MPORT_997_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_998_en & cosLUT_MPORT_998_mask) begin
      cosLUT[cosLUT_MPORT_998_addr] <= cosLUT_MPORT_998_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_999_en & cosLUT_MPORT_999_mask) begin
      cosLUT[cosLUT_MPORT_999_addr] <= cosLUT_MPORT_999_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1000_en & cosLUT_MPORT_1000_mask) begin
      cosLUT[cosLUT_MPORT_1000_addr] <= cosLUT_MPORT_1000_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1001_en & cosLUT_MPORT_1001_mask) begin
      cosLUT[cosLUT_MPORT_1001_addr] <= cosLUT_MPORT_1001_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1002_en & cosLUT_MPORT_1002_mask) begin
      cosLUT[cosLUT_MPORT_1002_addr] <= cosLUT_MPORT_1002_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1003_en & cosLUT_MPORT_1003_mask) begin
      cosLUT[cosLUT_MPORT_1003_addr] <= cosLUT_MPORT_1003_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1004_en & cosLUT_MPORT_1004_mask) begin
      cosLUT[cosLUT_MPORT_1004_addr] <= cosLUT_MPORT_1004_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1005_en & cosLUT_MPORT_1005_mask) begin
      cosLUT[cosLUT_MPORT_1005_addr] <= cosLUT_MPORT_1005_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1006_en & cosLUT_MPORT_1006_mask) begin
      cosLUT[cosLUT_MPORT_1006_addr] <= cosLUT_MPORT_1006_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1007_en & cosLUT_MPORT_1007_mask) begin
      cosLUT[cosLUT_MPORT_1007_addr] <= cosLUT_MPORT_1007_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1008_en & cosLUT_MPORT_1008_mask) begin
      cosLUT[cosLUT_MPORT_1008_addr] <= cosLUT_MPORT_1008_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1009_en & cosLUT_MPORT_1009_mask) begin
      cosLUT[cosLUT_MPORT_1009_addr] <= cosLUT_MPORT_1009_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1010_en & cosLUT_MPORT_1010_mask) begin
      cosLUT[cosLUT_MPORT_1010_addr] <= cosLUT_MPORT_1010_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1011_en & cosLUT_MPORT_1011_mask) begin
      cosLUT[cosLUT_MPORT_1011_addr] <= cosLUT_MPORT_1011_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1012_en & cosLUT_MPORT_1012_mask) begin
      cosLUT[cosLUT_MPORT_1012_addr] <= cosLUT_MPORT_1012_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1013_en & cosLUT_MPORT_1013_mask) begin
      cosLUT[cosLUT_MPORT_1013_addr] <= cosLUT_MPORT_1013_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1014_en & cosLUT_MPORT_1014_mask) begin
      cosLUT[cosLUT_MPORT_1014_addr] <= cosLUT_MPORT_1014_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1015_en & cosLUT_MPORT_1015_mask) begin
      cosLUT[cosLUT_MPORT_1015_addr] <= cosLUT_MPORT_1015_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1016_en & cosLUT_MPORT_1016_mask) begin
      cosLUT[cosLUT_MPORT_1016_addr] <= cosLUT_MPORT_1016_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1017_en & cosLUT_MPORT_1017_mask) begin
      cosLUT[cosLUT_MPORT_1017_addr] <= cosLUT_MPORT_1017_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1018_en & cosLUT_MPORT_1018_mask) begin
      cosLUT[cosLUT_MPORT_1018_addr] <= cosLUT_MPORT_1018_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1019_en & cosLUT_MPORT_1019_mask) begin
      cosLUT[cosLUT_MPORT_1019_addr] <= cosLUT_MPORT_1019_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1020_en & cosLUT_MPORT_1020_mask) begin
      cosLUT[cosLUT_MPORT_1020_addr] <= cosLUT_MPORT_1020_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1021_en & cosLUT_MPORT_1021_mask) begin
      cosLUT[cosLUT_MPORT_1021_addr] <= cosLUT_MPORT_1021_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1022_en & cosLUT_MPORT_1022_mask) begin
      cosLUT[cosLUT_MPORT_1022_addr] <= cosLUT_MPORT_1022_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1023_en & cosLUT_MPORT_1023_mask) begin
      cosLUT[cosLUT_MPORT_1023_addr] <= cosLUT_MPORT_1023_data; // @[LUTbank2.scala 323:29]
    end
    if (cosLUT_MPORT_1024_en & cosLUT_MPORT_1024_mask) begin
      cosLUT[cosLUT_MPORT_1024_addr] <= cosLUT_MPORT_1024_data; // @[LUTbank2.scala 323:29]
    end
    cosLUT_io_cosOut_0_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_0_MPORT_addr_pipe_0 <= io_cosIndex_0[10:0];
    end
    cosLUT_io_sinOut_0_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_0_MPORT_addr_pipe_0 <= io_sinIndex_0[10:0];
    end
    cosLUT_io_cosOut_1_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_1_MPORT_addr_pipe_0 <= io_cosIndex_1[10:0];
    end
    cosLUT_io_sinOut_1_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_1_MPORT_addr_pipe_0 <= io_sinIndex_1[10:0];
    end
    cosLUT_io_cosOut_2_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_2_MPORT_addr_pipe_0 <= io_cosIndex_2[10:0];
    end
    cosLUT_io_sinOut_2_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_2_MPORT_addr_pipe_0 <= io_sinIndex_2[10:0];
    end
    cosLUT_io_cosOut_3_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_3_MPORT_addr_pipe_0 <= io_cosIndex_3[10:0];
    end
    cosLUT_io_sinOut_3_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_3_MPORT_addr_pipe_0 <= io_sinIndex_3[10:0];
    end
    cosLUT_io_cosOut_4_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_4_MPORT_addr_pipe_0 <= io_cosIndex_4[10:0];
    end
    cosLUT_io_sinOut_4_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_4_MPORT_addr_pipe_0 <= io_sinIndex_4[10:0];
    end
    cosLUT_io_cosOut_5_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_5_MPORT_addr_pipe_0 <= io_cosIndex_5[10:0];
    end
    cosLUT_io_sinOut_5_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_5_MPORT_addr_pipe_0 <= io_sinIndex_5[10:0];
    end
    cosLUT_io_cosOut_6_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_6_MPORT_addr_pipe_0 <= io_cosIndex_6[10:0];
    end
    cosLUT_io_sinOut_6_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_6_MPORT_addr_pipe_0 <= io_sinIndex_6[10:0];
    end
    cosLUT_io_cosOut_7_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_cosOut_7_MPORT_addr_pipe_0 <= io_cosIndex_7[10:0];
    end
    cosLUT_io_sinOut_7_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cosLUT_io_sinOut_7_MPORT_addr_pipe_0 <= io_sinIndex_7[10:0];
    end
    if (reset) begin // @[LUTbank2.scala 331:29]
      ENReg <= 1'h0; // @[LUTbank2.scala 331:29]
    end else begin
      ENReg <= io_EN; // @[LUTbank2.scala 335:11]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_0_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_0_0 <= io_x_0_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_0_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_0_1 <= io_x_0_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_1_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_1_0 <= io_x_1_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_1_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_1_1 <= io_x_1_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_2_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_2_0 <= io_x_2_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_2_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_2_1 <= io_x_2_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_3_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_3_0 <= io_x_3_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_3_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_3_1 <= io_x_3_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_4_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_4_0 <= io_x_4_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_4_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_4_1 <= io_x_4_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_5_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_5_0 <= io_x_5_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_5_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_5_1 <= io_x_5_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_6_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_6_0 <= io_x_6_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_6_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_6_1 <= io_x_6_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_7_0 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_7_0 <= io_x_7_0; // @[LUTbank2.scala 337:23]
    end
    if (reset) begin // @[LUTbank2.scala 332:29]
      xFWDReg_7_1 <= 32'h0; // @[LUTbank2.scala 332:29]
    end else begin
      xFWDReg_7_1 <= io_x_7_1; // @[LUTbank2.scala 338:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_0_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_0_0 <= io_sign_0_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_0_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_0_1 <= io_sign_0_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_1_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_1_0 <= io_sign_1_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_1_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_1_1 <= io_sign_1_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_2_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_2_0 <= io_sign_2_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_2_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_2_1 <= io_sign_2_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_3_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_3_0 <= io_sign_3_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_3_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_3_1 <= io_sign_3_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_4_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_4_0 <= io_sign_4_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_4_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_4_1 <= io_sign_4_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_5_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_5_0 <= io_sign_5_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_5_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_5_1 <= io_sign_5_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_6_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_6_0 <= io_sign_6_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_6_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_6_1 <= io_sign_6_1; // @[LUTbank2.scala 340:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_7_0 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_7_0 <= io_sign_7_0; // @[LUTbank2.scala 339:23]
    end
    if (reset) begin // @[LUTbank2.scala 333:29]
      signReg_7_1 <= 1'h0; // @[LUTbank2.scala 333:29]
    end else begin
      signReg_7_1 <= io_sign_7_1; // @[LUTbank2.scala 340:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_8 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_10 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_12 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_14 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_16 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1025; initvar = initvar+1)
    cosLUT[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  cosLUT_io_cosOut_0_MPORT_en_pipe_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  cosLUT_io_cosOut_0_MPORT_addr_pipe_0 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  cosLUT_io_sinOut_0_MPORT_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cosLUT_io_sinOut_0_MPORT_addr_pipe_0 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  cosLUT_io_cosOut_1_MPORT_en_pipe_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  cosLUT_io_cosOut_1_MPORT_addr_pipe_0 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  cosLUT_io_sinOut_1_MPORT_en_pipe_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  cosLUT_io_sinOut_1_MPORT_addr_pipe_0 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  cosLUT_io_cosOut_2_MPORT_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cosLUT_io_cosOut_2_MPORT_addr_pipe_0 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  cosLUT_io_sinOut_2_MPORT_en_pipe_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  cosLUT_io_sinOut_2_MPORT_addr_pipe_0 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  cosLUT_io_cosOut_3_MPORT_en_pipe_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  cosLUT_io_cosOut_3_MPORT_addr_pipe_0 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  cosLUT_io_sinOut_3_MPORT_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cosLUT_io_sinOut_3_MPORT_addr_pipe_0 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  cosLUT_io_cosOut_4_MPORT_en_pipe_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  cosLUT_io_cosOut_4_MPORT_addr_pipe_0 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  cosLUT_io_sinOut_4_MPORT_en_pipe_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  cosLUT_io_sinOut_4_MPORT_addr_pipe_0 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  cosLUT_io_cosOut_5_MPORT_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  cosLUT_io_cosOut_5_MPORT_addr_pipe_0 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  cosLUT_io_sinOut_5_MPORT_en_pipe_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  cosLUT_io_sinOut_5_MPORT_addr_pipe_0 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  cosLUT_io_cosOut_6_MPORT_en_pipe_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  cosLUT_io_cosOut_6_MPORT_addr_pipe_0 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  cosLUT_io_sinOut_6_MPORT_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  cosLUT_io_sinOut_6_MPORT_addr_pipe_0 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  cosLUT_io_cosOut_7_MPORT_en_pipe_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cosLUT_io_cosOut_7_MPORT_addr_pipe_0 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  cosLUT_io_sinOut_7_MPORT_en_pipe_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  cosLUT_io_sinOut_7_MPORT_addr_pipe_0 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  ENReg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  xFWDReg_0_0 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  xFWDReg_0_1 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  xFWDReg_1_0 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  xFWDReg_1_1 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  xFWDReg_2_0 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  xFWDReg_2_1 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  xFWDReg_3_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  xFWDReg_3_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  xFWDReg_4_0 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  xFWDReg_4_1 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  xFWDReg_5_0 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  xFWDReg_5_1 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  xFWDReg_6_0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  xFWDReg_6_1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  xFWDReg_7_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  xFWDReg_7_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  signReg_0_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  signReg_0_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  signReg_1_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  signReg_1_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  signReg_2_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  signReg_2_1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  signReg_3_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  signReg_3_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  signReg_4_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  signReg_4_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  signReg_5_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  signReg_5_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  signReg_6_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  signReg_6_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  signReg_7_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  signReg_7_1 = _RAND_81[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module encoder(
  input         clock,
  input         reset,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input         io_EN,
  input  [31:0] io_cosIn,
  input  [31:0] io_sinIn,
  input         io_cosSign,
  input         io_sinSign,
  output [31:0] io_cosOut,
  output [31:0] io_sinOut,
  output        io_ENout,
  output [31:0] io_xFWD_0,
  output [31:0] io_xFWD_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  ENReg; // @[sincosLUT2.scala 134:29]
  reg [31:0] x0FWD; // @[sincosLUT2.scala 135:29]
  reg [31:0] x1FWD; // @[sincosLUT2.scala 136:29]
  reg [31:0] cosSign; // @[sincosLUT2.scala 137:29]
  reg [31:0] sinSign; // @[sincosLUT2.scala 138:29]
  reg [31:0] cos; // @[sincosLUT2.scala 139:29]
  reg [31:0] sin; // @[sincosLUT2.scala 140:29]
  wire [31:0] _GEN_0 = {{31'd0}, cos[31]}; // @[sincosLUT2.scala 150:31]
  wire [31:0] _io_cosOut_T_1 = cosSign ^ _GEN_0; // @[sincosLUT2.scala 150:31]
  wire [62:0] _io_cosOut_T_3 = {_io_cosOut_T_1,cos[30:0]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_1 = {{31'd0}, sin[31]}; // @[sincosLUT2.scala 151:31]
  wire [31:0] _io_sinOut_T_1 = sinSign ^ _GEN_1; // @[sincosLUT2.scala 151:31]
  wire [62:0] _io_sinOut_T_3 = {_io_sinOut_T_1,sin[30:0]}; // @[Cat.scala 33:92]
  assign io_cosOut = _io_cosOut_T_3[31:0]; // @[sincosLUT2.scala 150:16]
  assign io_sinOut = _io_sinOut_T_3[31:0]; // @[sincosLUT2.scala 151:16]
  assign io_ENout = ENReg; // @[sincosLUT2.scala 152:16]
  assign io_xFWD_0 = x0FWD; // @[sincosLUT2.scala 153:16]
  assign io_xFWD_1 = x1FWD; // @[sincosLUT2.scala 154:16]
  always @(posedge clock) begin
    if (reset) begin // @[sincosLUT2.scala 134:29]
      ENReg <= 1'h0; // @[sincosLUT2.scala 134:29]
    end else begin
      ENReg <= io_EN; // @[sincosLUT2.scala 142:13]
    end
    if (reset) begin // @[sincosLUT2.scala 135:29]
      x0FWD <= 32'h0; // @[sincosLUT2.scala 135:29]
    end else begin
      x0FWD <= io_x_0; // @[sincosLUT2.scala 143:13]
    end
    if (reset) begin // @[sincosLUT2.scala 136:29]
      x1FWD <= 32'h0; // @[sincosLUT2.scala 136:29]
    end else begin
      x1FWD <= io_x_1; // @[sincosLUT2.scala 144:13]
    end
    if (reset) begin // @[sincosLUT2.scala 137:29]
      cosSign <= 32'h0; // @[sincosLUT2.scala 137:29]
    end else begin
      cosSign <= {{31'd0}, io_cosSign}; // @[sincosLUT2.scala 145:13]
    end
    if (reset) begin // @[sincosLUT2.scala 138:29]
      sinSign <= 32'h0; // @[sincosLUT2.scala 138:29]
    end else begin
      sinSign <= {{31'd0}, io_sinSign}; // @[sincosLUT2.scala 146:13]
    end
    if (reset) begin // @[sincosLUT2.scala 139:29]
      cos <= 32'h0; // @[sincosLUT2.scala 139:29]
    end else begin
      cos <= io_cosIn; // @[sincosLUT2.scala 147:13]
    end
    if (reset) begin // @[sincosLUT2.scala 140:29]
      sin <= 32'h0; // @[sincosLUT2.scala 140:29]
    end else begin
      sin <= io_sinIn; // @[sincosLUT2.scala 148:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ENReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  x0FWD = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x1FWD = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cosSign = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  sinSign = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cos = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  sin = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multiPortSinCosModuleV2(
  input         clock,
  input         reset,
  input  [31:0] io_x_0_0,
  input  [31:0] io_x_0_1,
  input  [31:0] io_x_1_0,
  input  [31:0] io_x_1_1,
  input  [31:0] io_x_2_0,
  input  [31:0] io_x_2_1,
  input  [31:0] io_x_3_0,
  input  [31:0] io_x_3_1,
  input  [31:0] io_x_4_0,
  input  [31:0] io_x_4_1,
  input  [31:0] io_x_5_0,
  input  [31:0] io_x_5_1,
  input  [31:0] io_x_6_0,
  input  [31:0] io_x_6_1,
  input  [31:0] io_x_7_0,
  input  [31:0] io_x_7_1,
  input         io_EN,
  input  [31:0] io_angle_0,
  input  [31:0] io_angle_1,
  input  [31:0] io_angle_2,
  input  [31:0] io_angle_3,
  input  [31:0] io_angle_4,
  input  [31:0] io_angle_5,
  input  [31:0] io_angle_6,
  input  [31:0] io_angle_7,
  output [31:0] io_sinOut_0,
  output [31:0] io_sinOut_1,
  output [31:0] io_sinOut_2,
  output [31:0] io_sinOut_3,
  output [31:0] io_sinOut_4,
  output [31:0] io_sinOut_5,
  output [31:0] io_sinOut_6,
  output [31:0] io_sinOut_7,
  output [31:0] io_cosOut_0,
  output [31:0] io_cosOut_1,
  output [31:0] io_cosOut_2,
  output [31:0] io_cosOut_3,
  output [31:0] io_cosOut_4,
  output [31:0] io_cosOut_5,
  output [31:0] io_cosOut_6,
  output [31:0] io_cosOut_7,
  output        io_ENout,
  output [31:0] io_xFWD_0_0,
  output [31:0] io_xFWD_0_1,
  output [31:0] io_xFWD_1_0,
  output [31:0] io_xFWD_1_1,
  output [31:0] io_xFWD_2_0,
  output [31:0] io_xFWD_2_1,
  output [31:0] io_xFWD_3_0,
  output [31:0] io_xFWD_3_1,
  output [31:0] io_xFWD_4_0,
  output [31:0] io_xFWD_4_1,
  output [31:0] io_xFWD_5_0,
  output [31:0] io_xFWD_5_1,
  output [31:0] io_xFWD_6_0,
  output [31:0] io_xFWD_6_1,
  output [31:0] io_xFWD_7_0,
  output [31:0] io_xFWD_7_1
);
  wire  dualPortIndexCalculatorV2_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_1_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_1_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_2_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_2_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_3_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_3_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_4_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_4_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_5_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_5_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_6_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_6_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_clock; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_reset; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_x_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_x_1; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_io_EN; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_angle; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_cosIndex; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_sinIndex; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_io_cosSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_io_sinSign; // @[sincosLUT3.scala 67:15]
  wire  dualPortIndexCalculatorV2_7_io_ENout; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_xFWD_0; // @[sincosLUT3.scala 67:15]
  wire [31:0] dualPortIndexCalculatorV2_7_io_xFWD_1; // @[sincosLUT3.scala 67:15]
  wire  lutModule_clock; // @[sincosLUT3.scala 69:27]
  wire  lutModule_reset; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_EN; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_0_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_0_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_1_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_1_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_2_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_2_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_3_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_3_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_4_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_4_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_5_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_5_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_6_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_6_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_7_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_x_7_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_2; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_3; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_4; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_5; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_6; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosIndex_7; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_2; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_3; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_4; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_5; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_6; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinIndex_7; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_0_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_0_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_1_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_1_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_2_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_2_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_3_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_3_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_4_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_4_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_5_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_5_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_6_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_6_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_7_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_sign_7_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_2; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_3; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_4; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_5; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_6; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_sinOut_7; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_2; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_3; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_4; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_5; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_6; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_cosOut_7; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_ENout; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_0_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_0_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_1_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_1_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_2_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_2_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_3_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_3_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_4_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_4_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_5_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_5_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_6_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_6_1; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_7_0; // @[sincosLUT3.scala 69:27]
  wire [31:0] lutModule_io_xFWD_7_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_0_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_0_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_1_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_1_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_2_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_2_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_3_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_3_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_4_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_4_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_5_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_5_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_6_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_6_1; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_7_0; // @[sincosLUT3.scala 69:27]
  wire  lutModule_io_signFWD_7_1; // @[sincosLUT3.scala 69:27]
  wire  encoder_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_1_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_1_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_2_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_2_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_3_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_3_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_4_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_4_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_5_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_5_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_6_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_6_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_clock; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_reset; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_x_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_x_1; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_io_EN; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_cosIn; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_sinIn; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_io_cosSign; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_io_sinSign; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_cosOut; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_sinOut; // @[sincosLUT3.scala 71:15]
  wire  encoder_7_io_ENout; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_xFWD_0; // @[sincosLUT3.scala 71:15]
  wire [31:0] encoder_7_io_xFWD_1; // @[sincosLUT3.scala 71:15]
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_clock),
    .reset(dualPortIndexCalculatorV2_reset),
    .io_x_0(dualPortIndexCalculatorV2_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_io_EN),
    .io_angle(dualPortIndexCalculatorV2_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_1 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_1_clock),
    .reset(dualPortIndexCalculatorV2_1_reset),
    .io_x_0(dualPortIndexCalculatorV2_1_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_1_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_1_io_EN),
    .io_angle(dualPortIndexCalculatorV2_1_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_1_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_1_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_1_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_1_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_1_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_1_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_1_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_2 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_2_clock),
    .reset(dualPortIndexCalculatorV2_2_reset),
    .io_x_0(dualPortIndexCalculatorV2_2_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_2_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_2_io_EN),
    .io_angle(dualPortIndexCalculatorV2_2_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_2_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_2_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_2_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_2_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_2_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_2_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_2_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_3 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_3_clock),
    .reset(dualPortIndexCalculatorV2_3_reset),
    .io_x_0(dualPortIndexCalculatorV2_3_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_3_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_3_io_EN),
    .io_angle(dualPortIndexCalculatorV2_3_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_3_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_3_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_3_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_3_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_3_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_3_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_3_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_4 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_4_clock),
    .reset(dualPortIndexCalculatorV2_4_reset),
    .io_x_0(dualPortIndexCalculatorV2_4_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_4_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_4_io_EN),
    .io_angle(dualPortIndexCalculatorV2_4_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_4_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_4_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_4_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_4_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_4_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_4_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_4_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_5 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_5_clock),
    .reset(dualPortIndexCalculatorV2_5_reset),
    .io_x_0(dualPortIndexCalculatorV2_5_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_5_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_5_io_EN),
    .io_angle(dualPortIndexCalculatorV2_5_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_5_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_5_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_5_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_5_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_5_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_5_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_5_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_6 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_6_clock),
    .reset(dualPortIndexCalculatorV2_6_reset),
    .io_x_0(dualPortIndexCalculatorV2_6_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_6_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_6_io_EN),
    .io_angle(dualPortIndexCalculatorV2_6_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_6_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_6_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_6_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_6_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_6_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_6_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_6_io_xFWD_1)
  );
  dualPortIndexCalculatorV2 dualPortIndexCalculatorV2_7 ( // @[sincosLUT3.scala 67:15]
    .clock(dualPortIndexCalculatorV2_7_clock),
    .reset(dualPortIndexCalculatorV2_7_reset),
    .io_x_0(dualPortIndexCalculatorV2_7_io_x_0),
    .io_x_1(dualPortIndexCalculatorV2_7_io_x_1),
    .io_EN(dualPortIndexCalculatorV2_7_io_EN),
    .io_angle(dualPortIndexCalculatorV2_7_io_angle),
    .io_cosIndex(dualPortIndexCalculatorV2_7_io_cosIndex),
    .io_sinIndex(dualPortIndexCalculatorV2_7_io_sinIndex),
    .io_cosSign(dualPortIndexCalculatorV2_7_io_cosSign),
    .io_sinSign(dualPortIndexCalculatorV2_7_io_sinSign),
    .io_ENout(dualPortIndexCalculatorV2_7_io_ENout),
    .io_xFWD_0(dualPortIndexCalculatorV2_7_io_xFWD_0),
    .io_xFWD_1(dualPortIndexCalculatorV2_7_io_xFWD_1)
  );
  multiPortCOSlut lutModule ( // @[sincosLUT3.scala 69:27]
    .clock(lutModule_clock),
    .reset(lutModule_reset),
    .io_EN(lutModule_io_EN),
    .io_x_0_0(lutModule_io_x_0_0),
    .io_x_0_1(lutModule_io_x_0_1),
    .io_x_1_0(lutModule_io_x_1_0),
    .io_x_1_1(lutModule_io_x_1_1),
    .io_x_2_0(lutModule_io_x_2_0),
    .io_x_2_1(lutModule_io_x_2_1),
    .io_x_3_0(lutModule_io_x_3_0),
    .io_x_3_1(lutModule_io_x_3_1),
    .io_x_4_0(lutModule_io_x_4_0),
    .io_x_4_1(lutModule_io_x_4_1),
    .io_x_5_0(lutModule_io_x_5_0),
    .io_x_5_1(lutModule_io_x_5_1),
    .io_x_6_0(lutModule_io_x_6_0),
    .io_x_6_1(lutModule_io_x_6_1),
    .io_x_7_0(lutModule_io_x_7_0),
    .io_x_7_1(lutModule_io_x_7_1),
    .io_cosIndex_0(lutModule_io_cosIndex_0),
    .io_cosIndex_1(lutModule_io_cosIndex_1),
    .io_cosIndex_2(lutModule_io_cosIndex_2),
    .io_cosIndex_3(lutModule_io_cosIndex_3),
    .io_cosIndex_4(lutModule_io_cosIndex_4),
    .io_cosIndex_5(lutModule_io_cosIndex_5),
    .io_cosIndex_6(lutModule_io_cosIndex_6),
    .io_cosIndex_7(lutModule_io_cosIndex_7),
    .io_sinIndex_0(lutModule_io_sinIndex_0),
    .io_sinIndex_1(lutModule_io_sinIndex_1),
    .io_sinIndex_2(lutModule_io_sinIndex_2),
    .io_sinIndex_3(lutModule_io_sinIndex_3),
    .io_sinIndex_4(lutModule_io_sinIndex_4),
    .io_sinIndex_5(lutModule_io_sinIndex_5),
    .io_sinIndex_6(lutModule_io_sinIndex_6),
    .io_sinIndex_7(lutModule_io_sinIndex_7),
    .io_sign_0_0(lutModule_io_sign_0_0),
    .io_sign_0_1(lutModule_io_sign_0_1),
    .io_sign_1_0(lutModule_io_sign_1_0),
    .io_sign_1_1(lutModule_io_sign_1_1),
    .io_sign_2_0(lutModule_io_sign_2_0),
    .io_sign_2_1(lutModule_io_sign_2_1),
    .io_sign_3_0(lutModule_io_sign_3_0),
    .io_sign_3_1(lutModule_io_sign_3_1),
    .io_sign_4_0(lutModule_io_sign_4_0),
    .io_sign_4_1(lutModule_io_sign_4_1),
    .io_sign_5_0(lutModule_io_sign_5_0),
    .io_sign_5_1(lutModule_io_sign_5_1),
    .io_sign_6_0(lutModule_io_sign_6_0),
    .io_sign_6_1(lutModule_io_sign_6_1),
    .io_sign_7_0(lutModule_io_sign_7_0),
    .io_sign_7_1(lutModule_io_sign_7_1),
    .io_sinOut_0(lutModule_io_sinOut_0),
    .io_sinOut_1(lutModule_io_sinOut_1),
    .io_sinOut_2(lutModule_io_sinOut_2),
    .io_sinOut_3(lutModule_io_sinOut_3),
    .io_sinOut_4(lutModule_io_sinOut_4),
    .io_sinOut_5(lutModule_io_sinOut_5),
    .io_sinOut_6(lutModule_io_sinOut_6),
    .io_sinOut_7(lutModule_io_sinOut_7),
    .io_cosOut_0(lutModule_io_cosOut_0),
    .io_cosOut_1(lutModule_io_cosOut_1),
    .io_cosOut_2(lutModule_io_cosOut_2),
    .io_cosOut_3(lutModule_io_cosOut_3),
    .io_cosOut_4(lutModule_io_cosOut_4),
    .io_cosOut_5(lutModule_io_cosOut_5),
    .io_cosOut_6(lutModule_io_cosOut_6),
    .io_cosOut_7(lutModule_io_cosOut_7),
    .io_ENout(lutModule_io_ENout),
    .io_xFWD_0_0(lutModule_io_xFWD_0_0),
    .io_xFWD_0_1(lutModule_io_xFWD_0_1),
    .io_xFWD_1_0(lutModule_io_xFWD_1_0),
    .io_xFWD_1_1(lutModule_io_xFWD_1_1),
    .io_xFWD_2_0(lutModule_io_xFWD_2_0),
    .io_xFWD_2_1(lutModule_io_xFWD_2_1),
    .io_xFWD_3_0(lutModule_io_xFWD_3_0),
    .io_xFWD_3_1(lutModule_io_xFWD_3_1),
    .io_xFWD_4_0(lutModule_io_xFWD_4_0),
    .io_xFWD_4_1(lutModule_io_xFWD_4_1),
    .io_xFWD_5_0(lutModule_io_xFWD_5_0),
    .io_xFWD_5_1(lutModule_io_xFWD_5_1),
    .io_xFWD_6_0(lutModule_io_xFWD_6_0),
    .io_xFWD_6_1(lutModule_io_xFWD_6_1),
    .io_xFWD_7_0(lutModule_io_xFWD_7_0),
    .io_xFWD_7_1(lutModule_io_xFWD_7_1),
    .io_signFWD_0_0(lutModule_io_signFWD_0_0),
    .io_signFWD_0_1(lutModule_io_signFWD_0_1),
    .io_signFWD_1_0(lutModule_io_signFWD_1_0),
    .io_signFWD_1_1(lutModule_io_signFWD_1_1),
    .io_signFWD_2_0(lutModule_io_signFWD_2_0),
    .io_signFWD_2_1(lutModule_io_signFWD_2_1),
    .io_signFWD_3_0(lutModule_io_signFWD_3_0),
    .io_signFWD_3_1(lutModule_io_signFWD_3_1),
    .io_signFWD_4_0(lutModule_io_signFWD_4_0),
    .io_signFWD_4_1(lutModule_io_signFWD_4_1),
    .io_signFWD_5_0(lutModule_io_signFWD_5_0),
    .io_signFWD_5_1(lutModule_io_signFWD_5_1),
    .io_signFWD_6_0(lutModule_io_signFWD_6_0),
    .io_signFWD_6_1(lutModule_io_signFWD_6_1),
    .io_signFWD_7_0(lutModule_io_signFWD_7_0),
    .io_signFWD_7_1(lutModule_io_signFWD_7_1)
  );
  encoder encoder ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_clock),
    .reset(encoder_reset),
    .io_x_0(encoder_io_x_0),
    .io_x_1(encoder_io_x_1),
    .io_EN(encoder_io_EN),
    .io_cosIn(encoder_io_cosIn),
    .io_sinIn(encoder_io_sinIn),
    .io_cosSign(encoder_io_cosSign),
    .io_sinSign(encoder_io_sinSign),
    .io_cosOut(encoder_io_cosOut),
    .io_sinOut(encoder_io_sinOut),
    .io_ENout(encoder_io_ENout),
    .io_xFWD_0(encoder_io_xFWD_0),
    .io_xFWD_1(encoder_io_xFWD_1)
  );
  encoder encoder_1 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_1_clock),
    .reset(encoder_1_reset),
    .io_x_0(encoder_1_io_x_0),
    .io_x_1(encoder_1_io_x_1),
    .io_EN(encoder_1_io_EN),
    .io_cosIn(encoder_1_io_cosIn),
    .io_sinIn(encoder_1_io_sinIn),
    .io_cosSign(encoder_1_io_cosSign),
    .io_sinSign(encoder_1_io_sinSign),
    .io_cosOut(encoder_1_io_cosOut),
    .io_sinOut(encoder_1_io_sinOut),
    .io_ENout(encoder_1_io_ENout),
    .io_xFWD_0(encoder_1_io_xFWD_0),
    .io_xFWD_1(encoder_1_io_xFWD_1)
  );
  encoder encoder_2 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_2_clock),
    .reset(encoder_2_reset),
    .io_x_0(encoder_2_io_x_0),
    .io_x_1(encoder_2_io_x_1),
    .io_EN(encoder_2_io_EN),
    .io_cosIn(encoder_2_io_cosIn),
    .io_sinIn(encoder_2_io_sinIn),
    .io_cosSign(encoder_2_io_cosSign),
    .io_sinSign(encoder_2_io_sinSign),
    .io_cosOut(encoder_2_io_cosOut),
    .io_sinOut(encoder_2_io_sinOut),
    .io_ENout(encoder_2_io_ENout),
    .io_xFWD_0(encoder_2_io_xFWD_0),
    .io_xFWD_1(encoder_2_io_xFWD_1)
  );
  encoder encoder_3 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_3_clock),
    .reset(encoder_3_reset),
    .io_x_0(encoder_3_io_x_0),
    .io_x_1(encoder_3_io_x_1),
    .io_EN(encoder_3_io_EN),
    .io_cosIn(encoder_3_io_cosIn),
    .io_sinIn(encoder_3_io_sinIn),
    .io_cosSign(encoder_3_io_cosSign),
    .io_sinSign(encoder_3_io_sinSign),
    .io_cosOut(encoder_3_io_cosOut),
    .io_sinOut(encoder_3_io_sinOut),
    .io_ENout(encoder_3_io_ENout),
    .io_xFWD_0(encoder_3_io_xFWD_0),
    .io_xFWD_1(encoder_3_io_xFWD_1)
  );
  encoder encoder_4 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_4_clock),
    .reset(encoder_4_reset),
    .io_x_0(encoder_4_io_x_0),
    .io_x_1(encoder_4_io_x_1),
    .io_EN(encoder_4_io_EN),
    .io_cosIn(encoder_4_io_cosIn),
    .io_sinIn(encoder_4_io_sinIn),
    .io_cosSign(encoder_4_io_cosSign),
    .io_sinSign(encoder_4_io_sinSign),
    .io_cosOut(encoder_4_io_cosOut),
    .io_sinOut(encoder_4_io_sinOut),
    .io_ENout(encoder_4_io_ENout),
    .io_xFWD_0(encoder_4_io_xFWD_0),
    .io_xFWD_1(encoder_4_io_xFWD_1)
  );
  encoder encoder_5 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_5_clock),
    .reset(encoder_5_reset),
    .io_x_0(encoder_5_io_x_0),
    .io_x_1(encoder_5_io_x_1),
    .io_EN(encoder_5_io_EN),
    .io_cosIn(encoder_5_io_cosIn),
    .io_sinIn(encoder_5_io_sinIn),
    .io_cosSign(encoder_5_io_cosSign),
    .io_sinSign(encoder_5_io_sinSign),
    .io_cosOut(encoder_5_io_cosOut),
    .io_sinOut(encoder_5_io_sinOut),
    .io_ENout(encoder_5_io_ENout),
    .io_xFWD_0(encoder_5_io_xFWD_0),
    .io_xFWD_1(encoder_5_io_xFWD_1)
  );
  encoder encoder_6 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_6_clock),
    .reset(encoder_6_reset),
    .io_x_0(encoder_6_io_x_0),
    .io_x_1(encoder_6_io_x_1),
    .io_EN(encoder_6_io_EN),
    .io_cosIn(encoder_6_io_cosIn),
    .io_sinIn(encoder_6_io_sinIn),
    .io_cosSign(encoder_6_io_cosSign),
    .io_sinSign(encoder_6_io_sinSign),
    .io_cosOut(encoder_6_io_cosOut),
    .io_sinOut(encoder_6_io_sinOut),
    .io_ENout(encoder_6_io_ENout),
    .io_xFWD_0(encoder_6_io_xFWD_0),
    .io_xFWD_1(encoder_6_io_xFWD_1)
  );
  encoder encoder_7 ( // @[sincosLUT3.scala 71:15]
    .clock(encoder_7_clock),
    .reset(encoder_7_reset),
    .io_x_0(encoder_7_io_x_0),
    .io_x_1(encoder_7_io_x_1),
    .io_EN(encoder_7_io_EN),
    .io_cosIn(encoder_7_io_cosIn),
    .io_sinIn(encoder_7_io_sinIn),
    .io_cosSign(encoder_7_io_cosSign),
    .io_sinSign(encoder_7_io_sinSign),
    .io_cosOut(encoder_7_io_cosOut),
    .io_sinOut(encoder_7_io_sinOut),
    .io_ENout(encoder_7_io_ENout),
    .io_xFWD_0(encoder_7_io_xFWD_0),
    .io_xFWD_1(encoder_7_io_xFWD_1)
  );
  assign io_sinOut_0 = encoder_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_1 = encoder_1_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_2 = encoder_2_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_3 = encoder_3_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_4 = encoder_4_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_5 = encoder_5_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_6 = encoder_6_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_sinOut_7 = encoder_7_io_sinOut; // @[sincosLUT3.scala 110:23]
  assign io_cosOut_0 = encoder_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_1 = encoder_1_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_2 = encoder_2_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_3 = encoder_3_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_4 = encoder_4_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_5 = encoder_5_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_6 = encoder_6_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_cosOut_7 = encoder_7_io_cosOut; // @[sincosLUT3.scala 109:23]
  assign io_ENout = encoder_io_ENout; // @[sincosLUT3.scala 105:23]
  assign io_xFWD_0_0 = encoder_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_0_1 = encoder_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_1_0 = encoder_1_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_1_1 = encoder_1_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_2_0 = encoder_2_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_2_1 = encoder_2_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_3_0 = encoder_3_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_3_1 = encoder_3_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_4_0 = encoder_4_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_4_1 = encoder_4_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_5_0 = encoder_5_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_5_1 = encoder_5_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_6_0 = encoder_6_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_6_1 = encoder_6_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign io_xFWD_7_0 = encoder_7_io_xFWD_0; // @[sincosLUT3.scala 107:23]
  assign io_xFWD_7_1 = encoder_7_io_xFWD_1; // @[sincosLUT3.scala 108:23]
  assign dualPortIndexCalculatorV2_clock = clock;
  assign dualPortIndexCalculatorV2_reset = reset;
  assign dualPortIndexCalculatorV2_io_x_0 = io_x_0_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_io_x_1 = io_x_0_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_io_angle = io_angle_0; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_1_clock = clock;
  assign dualPortIndexCalculatorV2_1_reset = reset;
  assign dualPortIndexCalculatorV2_1_io_x_0 = io_x_1_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_1_io_x_1 = io_x_1_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_1_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_1_io_angle = io_angle_1; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_2_clock = clock;
  assign dualPortIndexCalculatorV2_2_reset = reset;
  assign dualPortIndexCalculatorV2_2_io_x_0 = io_x_2_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_2_io_x_1 = io_x_2_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_2_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_2_io_angle = io_angle_2; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_3_clock = clock;
  assign dualPortIndexCalculatorV2_3_reset = reset;
  assign dualPortIndexCalculatorV2_3_io_x_0 = io_x_3_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_3_io_x_1 = io_x_3_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_3_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_3_io_angle = io_angle_3; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_4_clock = clock;
  assign dualPortIndexCalculatorV2_4_reset = reset;
  assign dualPortIndexCalculatorV2_4_io_x_0 = io_x_4_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_4_io_x_1 = io_x_4_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_4_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_4_io_angle = io_angle_4; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_5_clock = clock;
  assign dualPortIndexCalculatorV2_5_reset = reset;
  assign dualPortIndexCalculatorV2_5_io_x_0 = io_x_5_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_5_io_x_1 = io_x_5_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_5_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_5_io_angle = io_angle_5; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_6_clock = clock;
  assign dualPortIndexCalculatorV2_6_reset = reset;
  assign dualPortIndexCalculatorV2_6_io_x_0 = io_x_6_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_6_io_x_1 = io_x_6_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_6_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_6_io_angle = io_angle_6; // @[sincosLUT3.scala 79:37]
  assign dualPortIndexCalculatorV2_7_clock = clock;
  assign dualPortIndexCalculatorV2_7_reset = reset;
  assign dualPortIndexCalculatorV2_7_io_x_0 = io_x_7_0; // @[sincosLUT3.scala 77:37]
  assign dualPortIndexCalculatorV2_7_io_x_1 = io_x_7_1; // @[sincosLUT3.scala 78:37]
  assign dualPortIndexCalculatorV2_7_io_EN = io_EN; // @[sincosLUT3.scala 76:37]
  assign dualPortIndexCalculatorV2_7_io_angle = io_angle_7; // @[sincosLUT3.scala 79:37]
  assign lutModule_clock = clock;
  assign lutModule_reset = reset;
  assign lutModule_io_EN = dualPortIndexCalculatorV2_io_ENout; // @[sincosLUT3.scala 83:37]
  assign lutModule_io_x_0_0 = dualPortIndexCalculatorV2_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_0_1 = dualPortIndexCalculatorV2_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_1_0 = dualPortIndexCalculatorV2_1_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_1_1 = dualPortIndexCalculatorV2_1_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_2_0 = dualPortIndexCalculatorV2_2_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_2_1 = dualPortIndexCalculatorV2_2_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_3_0 = dualPortIndexCalculatorV2_3_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_3_1 = dualPortIndexCalculatorV2_3_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_4_0 = dualPortIndexCalculatorV2_4_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_4_1 = dualPortIndexCalculatorV2_4_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_5_0 = dualPortIndexCalculatorV2_5_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_5_1 = dualPortIndexCalculatorV2_5_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_6_0 = dualPortIndexCalculatorV2_6_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_6_1 = dualPortIndexCalculatorV2_6_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_x_7_0 = dualPortIndexCalculatorV2_7_io_xFWD_0; // @[sincosLUT3.scala 85:37]
  assign lutModule_io_x_7_1 = dualPortIndexCalculatorV2_7_io_xFWD_1; // @[sincosLUT3.scala 86:37]
  assign lutModule_io_cosIndex_0 = dualPortIndexCalculatorV2_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_1 = dualPortIndexCalculatorV2_1_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_2 = dualPortIndexCalculatorV2_2_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_3 = dualPortIndexCalculatorV2_3_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_4 = dualPortIndexCalculatorV2_4_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_5 = dualPortIndexCalculatorV2_5_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_6 = dualPortIndexCalculatorV2_6_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_cosIndex_7 = dualPortIndexCalculatorV2_7_io_cosIndex; // @[sincosLUT3.scala 87:37]
  assign lutModule_io_sinIndex_0 = dualPortIndexCalculatorV2_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_1 = dualPortIndexCalculatorV2_1_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_2 = dualPortIndexCalculatorV2_2_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_3 = dualPortIndexCalculatorV2_3_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_4 = dualPortIndexCalculatorV2_4_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_5 = dualPortIndexCalculatorV2_5_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_6 = dualPortIndexCalculatorV2_6_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sinIndex_7 = dualPortIndexCalculatorV2_7_io_sinIndex; // @[sincosLUT3.scala 88:37]
  assign lutModule_io_sign_0_0 = dualPortIndexCalculatorV2_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_0_1 = dualPortIndexCalculatorV2_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_1_0 = dualPortIndexCalculatorV2_1_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_1_1 = dualPortIndexCalculatorV2_1_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_2_0 = dualPortIndexCalculatorV2_2_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_2_1 = dualPortIndexCalculatorV2_2_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_3_0 = dualPortIndexCalculatorV2_3_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_3_1 = dualPortIndexCalculatorV2_3_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_4_0 = dualPortIndexCalculatorV2_4_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_4_1 = dualPortIndexCalculatorV2_4_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_5_0 = dualPortIndexCalculatorV2_5_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_5_1 = dualPortIndexCalculatorV2_5_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_6_0 = dualPortIndexCalculatorV2_6_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_6_1 = dualPortIndexCalculatorV2_6_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign lutModule_io_sign_7_0 = dualPortIndexCalculatorV2_7_io_cosSign; // @[sincosLUT3.scala 89:37]
  assign lutModule_io_sign_7_1 = dualPortIndexCalculatorV2_7_io_sinSign; // @[sincosLUT3.scala 90:37]
  assign encoder_clock = clock;
  assign encoder_reset = reset;
  assign encoder_io_x_0 = lutModule_io_xFWD_0_0; // @[sincosLUT3.scala 96:31]
  assign encoder_io_x_1 = lutModule_io_xFWD_0_1; // @[sincosLUT3.scala 97:31]
  assign encoder_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_io_cosIn = lutModule_io_cosOut_0; // @[sincosLUT3.scala 98:31]
  assign encoder_io_sinIn = lutModule_io_sinOut_0; // @[sincosLUT3.scala 99:31]
  assign encoder_io_cosSign = lutModule_io_signFWD_0_0; // @[sincosLUT3.scala 100:31]
  assign encoder_io_sinSign = lutModule_io_signFWD_0_1; // @[sincosLUT3.scala 101:31]
  assign encoder_1_clock = clock;
  assign encoder_1_reset = reset;
  assign encoder_1_io_x_0 = lutModule_io_xFWD_1_0; // @[sincosLUT3.scala 96:31]
  assign encoder_1_io_x_1 = lutModule_io_xFWD_1_1; // @[sincosLUT3.scala 97:31]
  assign encoder_1_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_1_io_cosIn = lutModule_io_cosOut_1; // @[sincosLUT3.scala 98:31]
  assign encoder_1_io_sinIn = lutModule_io_sinOut_1; // @[sincosLUT3.scala 99:31]
  assign encoder_1_io_cosSign = lutModule_io_signFWD_1_0; // @[sincosLUT3.scala 100:31]
  assign encoder_1_io_sinSign = lutModule_io_signFWD_1_1; // @[sincosLUT3.scala 101:31]
  assign encoder_2_clock = clock;
  assign encoder_2_reset = reset;
  assign encoder_2_io_x_0 = lutModule_io_xFWD_2_0; // @[sincosLUT3.scala 96:31]
  assign encoder_2_io_x_1 = lutModule_io_xFWD_2_1; // @[sincosLUT3.scala 97:31]
  assign encoder_2_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_2_io_cosIn = lutModule_io_cosOut_2; // @[sincosLUT3.scala 98:31]
  assign encoder_2_io_sinIn = lutModule_io_sinOut_2; // @[sincosLUT3.scala 99:31]
  assign encoder_2_io_cosSign = lutModule_io_signFWD_2_0; // @[sincosLUT3.scala 100:31]
  assign encoder_2_io_sinSign = lutModule_io_signFWD_2_1; // @[sincosLUT3.scala 101:31]
  assign encoder_3_clock = clock;
  assign encoder_3_reset = reset;
  assign encoder_3_io_x_0 = lutModule_io_xFWD_3_0; // @[sincosLUT3.scala 96:31]
  assign encoder_3_io_x_1 = lutModule_io_xFWD_3_1; // @[sincosLUT3.scala 97:31]
  assign encoder_3_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_3_io_cosIn = lutModule_io_cosOut_3; // @[sincosLUT3.scala 98:31]
  assign encoder_3_io_sinIn = lutModule_io_sinOut_3; // @[sincosLUT3.scala 99:31]
  assign encoder_3_io_cosSign = lutModule_io_signFWD_3_0; // @[sincosLUT3.scala 100:31]
  assign encoder_3_io_sinSign = lutModule_io_signFWD_3_1; // @[sincosLUT3.scala 101:31]
  assign encoder_4_clock = clock;
  assign encoder_4_reset = reset;
  assign encoder_4_io_x_0 = lutModule_io_xFWD_4_0; // @[sincosLUT3.scala 96:31]
  assign encoder_4_io_x_1 = lutModule_io_xFWD_4_1; // @[sincosLUT3.scala 97:31]
  assign encoder_4_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_4_io_cosIn = lutModule_io_cosOut_4; // @[sincosLUT3.scala 98:31]
  assign encoder_4_io_sinIn = lutModule_io_sinOut_4; // @[sincosLUT3.scala 99:31]
  assign encoder_4_io_cosSign = lutModule_io_signFWD_4_0; // @[sincosLUT3.scala 100:31]
  assign encoder_4_io_sinSign = lutModule_io_signFWD_4_1; // @[sincosLUT3.scala 101:31]
  assign encoder_5_clock = clock;
  assign encoder_5_reset = reset;
  assign encoder_5_io_x_0 = lutModule_io_xFWD_5_0; // @[sincosLUT3.scala 96:31]
  assign encoder_5_io_x_1 = lutModule_io_xFWD_5_1; // @[sincosLUT3.scala 97:31]
  assign encoder_5_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_5_io_cosIn = lutModule_io_cosOut_5; // @[sincosLUT3.scala 98:31]
  assign encoder_5_io_sinIn = lutModule_io_sinOut_5; // @[sincosLUT3.scala 99:31]
  assign encoder_5_io_cosSign = lutModule_io_signFWD_5_0; // @[sincosLUT3.scala 100:31]
  assign encoder_5_io_sinSign = lutModule_io_signFWD_5_1; // @[sincosLUT3.scala 101:31]
  assign encoder_6_clock = clock;
  assign encoder_6_reset = reset;
  assign encoder_6_io_x_0 = lutModule_io_xFWD_6_0; // @[sincosLUT3.scala 96:31]
  assign encoder_6_io_x_1 = lutModule_io_xFWD_6_1; // @[sincosLUT3.scala 97:31]
  assign encoder_6_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_6_io_cosIn = lutModule_io_cosOut_6; // @[sincosLUT3.scala 98:31]
  assign encoder_6_io_sinIn = lutModule_io_sinOut_6; // @[sincosLUT3.scala 99:31]
  assign encoder_6_io_cosSign = lutModule_io_signFWD_6_0; // @[sincosLUT3.scala 100:31]
  assign encoder_6_io_sinSign = lutModule_io_signFWD_6_1; // @[sincosLUT3.scala 101:31]
  assign encoder_7_clock = clock;
  assign encoder_7_reset = reset;
  assign encoder_7_io_x_0 = lutModule_io_xFWD_7_0; // @[sincosLUT3.scala 96:31]
  assign encoder_7_io_x_1 = lutModule_io_xFWD_7_1; // @[sincosLUT3.scala 97:31]
  assign encoder_7_io_EN = lutModule_io_ENout; // @[sincosLUT3.scala 95:31]
  assign encoder_7_io_cosIn = lutModule_io_cosOut_7; // @[sincosLUT3.scala 98:31]
  assign encoder_7_io_sinIn = lutModule_io_sinOut_7; // @[sincosLUT3.scala 99:31]
  assign encoder_7_io_cosSign = lutModule_io_signFWD_7_0; // @[sincosLUT3.scala 100:31]
  assign encoder_7_io_sinSign = lutModule_io_signFWD_7_1; // @[sincosLUT3.scala 101:31]
endmodule
module MulFullRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [47:0] io_rawOut_sig
);
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isZero | io_a_isZero & io_b_isInf; // @[MulRecFN.scala 58:60]
  wire [9:0] _common_sExpOut_T_2 = $signed(io_a_sExp) + $signed(io_b_sExp); // @[MulRecFN.scala 62:36]
  wire [49:0] _common_sigOut_T = io_a_sig * io_b_sig; // @[MulRecFN.scala 63:35]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[MulRecFN.scala 66:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[MulRecFN.scala 70:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[MulRecFN.scala 59:38]
  assign io_rawOut_isZero = io_a_isZero | io_b_isZero; // @[MulRecFN.scala 60:40]
  assign io_rawOut_sign = io_a_sign ^ io_b_sign; // @[MulRecFN.scala 61:36]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - 10'sh100; // @[MulRecFN.scala 62:48]
  assign io_rawOut_sig = _common_sigOut_T[47:0]; // @[MulRecFN.scala 63:46]
endmodule
module MulRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  mulFullRaw_io_a_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_a_sExp; // @[MulRecFN.scala 84:28]
  wire [24:0] mulFullRaw_io_a_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_b_sExp; // @[MulRecFN.scala 84:28]
  wire [24:0] mulFullRaw_io_b_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_invalidExc; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 84:28]
  wire [9:0] mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 84:28]
  wire [47:0] mulFullRaw_io_rawOut_sig; // @[MulRecFN.scala 84:28]
  wire  _io_rawOut_sig_T_2 = |mulFullRaw_io_rawOut_sig[21:0]; // @[MulRecFN.scala 93:55]
  MulFullRawFN mulFullRaw ( // @[MulRecFN.scala 84:28]
    .io_a_isNaN(mulFullRaw_io_a_isNaN),
    .io_a_isInf(mulFullRaw_io_a_isInf),
    .io_a_isZero(mulFullRaw_io_a_isZero),
    .io_a_sign(mulFullRaw_io_a_sign),
    .io_a_sExp(mulFullRaw_io_a_sExp),
    .io_a_sig(mulFullRaw_io_a_sig),
    .io_b_isNaN(mulFullRaw_io_b_isNaN),
    .io_b_isInf(mulFullRaw_io_b_isInf),
    .io_b_isZero(mulFullRaw_io_b_isZero),
    .io_b_sign(mulFullRaw_io_b_sign),
    .io_b_sExp(mulFullRaw_io_b_sExp),
    .io_b_sig(mulFullRaw_io_b_sig),
    .io_invalidExc(mulFullRaw_io_invalidExc),
    .io_rawOut_isNaN(mulFullRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(mulFullRaw_io_rawOut_isInf),
    .io_rawOut_isZero(mulFullRaw_io_rawOut_isZero),
    .io_rawOut_sign(mulFullRaw_io_rawOut_sign),
    .io_rawOut_sExp(mulFullRaw_io_rawOut_sExp),
    .io_rawOut_sig(mulFullRaw_io_rawOut_sig)
  );
  assign io_invalidExc = mulFullRaw_io_invalidExc; // @[MulRecFN.scala 89:19]
  assign io_rawOut_isNaN = mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isInf = mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isZero = mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sign = mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sExp = mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sig = {mulFullRaw_io_rawOut_sig[47:22],_io_rawOut_sig_T_2}; // @[Cat.scala 33:92]
  assign mulFullRaw_io_a_isNaN = io_a_isNaN; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isInf = io_a_isInf; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isZero = io_a_isZero; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sign = io_a_sign; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sExp = io_a_sExp; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sig = io_a_sig; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_b_isNaN = io_b_isNaN; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isInf = io_b_isInf; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isZero = io_b_isZero; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sign = io_b_sign; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sExp = io_b_sExp; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sig = io_b_sig; // @[MulRecFN.scala 87:21]
endmodule
module RoundAnyRawFNToRecFN_ie8_is26_oe8_os24(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 120:57]
  wire [8:0] _roundMask_T_1 = ~io_in_sExp[8:0]; // @[primitives.scala 52:21]
  wire  roundMask_msb = _roundMask_T_1[8]; // @[primitives.scala 58:25]
  wire [7:0] roundMask_lsbs = _roundMask_T_1[7:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_1 = roundMask_lsbs[7]; // @[primitives.scala 58:25]
  wire [6:0] roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[6]; // @[primitives.scala 58:25]
  wire [5:0] roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[primitives.scala 59:26]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> roundMask_lsbs_2; // @[primitives.scala 76:56]
  wire [15:0] _GEN_0 = {{8'd0}, roundMask_shift[57:50]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_7 = _GEN_0 & 16'hff; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_9 = {roundMask_shift[49:42], 8'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_11 = _roundMask_T_9 & 16'hff00; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_1 = {{4'd0}, _roundMask_T_12[15:4]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_17 = _GEN_1 & 16'hf0f; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_19 = {_roundMask_T_12[11:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_21 = _roundMask_T_19 & 16'hf0f0; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_2 = {{2'd0}, _roundMask_T_22[15:2]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_27 = _GEN_2 & 16'h3333; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_29 = {_roundMask_T_22[13:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_31 = _roundMask_T_29 & 16'hcccc; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 108:39]
  wire [15:0] _GEN_3 = {{1'd0}, _roundMask_T_32[15:1]}; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_37 = _GEN_3 & 16'h5555; // @[Bitwise.scala 108:31]
  wire [15:0] _roundMask_T_39 = {_roundMask_T_32[14:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [15:0] _roundMask_T_41 = _roundMask_T_39 & 16'haaaa; // @[Bitwise.scala 108:80]
  wire [15:0] _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 108:39]
  wire [21:0] _roundMask_T_59 = {_roundMask_T_42,roundMask_shift[58],roundMask_shift[59],roundMask_shift[60],
    roundMask_shift[61],roundMask_shift[62],roundMask_shift[63]}; // @[Cat.scala 33:92]
  wire [21:0] _roundMask_T_60 = ~_roundMask_T_59; // @[primitives.scala 73:32]
  wire [21:0] _roundMask_T_61 = roundMask_msb_2 ? 22'h0 : _roundMask_T_60; // @[primitives.scala 73:21]
  wire [21:0] _roundMask_T_62 = ~_roundMask_T_61; // @[primitives.scala 73:17]
  wire [24:0] _roundMask_T_63 = {_roundMask_T_62,3'h7}; // @[primitives.scala 68:58]
  wire [2:0] _roundMask_T_70 = {roundMask_shift[0],roundMask_shift[1],roundMask_shift[2]}; // @[Cat.scala 33:92]
  wire [2:0] _roundMask_T_71 = roundMask_msb_2 ? _roundMask_T_70 : 3'h0; // @[primitives.scala 62:24]
  wire [24:0] _roundMask_T_72 = roundMask_msb_1 ? _roundMask_T_63 : {{22'd0}, _roundMask_T_71}; // @[primitives.scala 67:24]
  wire [24:0] _roundMask_T_73 = roundMask_msb ? _roundMask_T_72 : 25'h0; // @[primitives.scala 62:24]
  wire [24:0] _GEN_4 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [24:0] _roundMask_T_74 = _roundMask_T_73 | _GEN_4; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [26:0] roundMask = {_roundMask_T_74,2'h3}; // @[RoundAnyRawFNToRecFN.scala 159:42]
  wire [27:0] _shiftedRoundMask_T = {1'h0,_roundMask_T_74,2'h3}; // @[RoundAnyRawFNToRecFN.scala 162:41]
  wire [26:0] shiftedRoundMask = _shiftedRoundMask_T[27:1]; // @[RoundAnyRawFNToRecFN.scala 162:53]
  wire [26:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:28]
  wire [26:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 163:46]
  wire [26:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 164:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 164:56]
  wire [26:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 165:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 165:62]
  wire [26:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 174:32]
  wire [25:0] _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 174:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 176:30]
  wire [25:0] _roundedSig_T_7 = roundPosBit & _roundedSig_T_4 ? roundMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 175:25]
  wire [25:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 175:21]
  wire [25:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 174:57]
  wire [26:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 180:32]
  wire [26:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 180:30]
  wire [25:0] _roundedSig_T_16 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 180:47]
  wire [25:0] roundedSig = roundPosBit ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 173:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 185:76]
  wire [9:0] _GEN_5 = {{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [10:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [8:0] common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 187:37]
  wire [22:0] common_fractOut = doShiftSigDown1 ? roundedSig[23:1] : roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:16]
  wire [3:0] _common_overflow_T = sRoundedExp[10:7]; // @[RoundAnyRawFNToRecFN.scala 196:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 196:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 200:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 235:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 237:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 238:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 248:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 250:22]
  wire [8:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 253:18]
  wire [8:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 253:14]
  wire [8:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 252:24]
  wire [8:0] _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 265:18]
  wire [8:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 265:14]
  wire [8:0] _expOut_T_13 = _expOut_T_3 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 264:17]
  wire [8:0] _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 277:16]
  wire [8:0] _expOut_T_19 = _expOut_T_13 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 276:15]
  wire [8:0] _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 278:16]
  wire [8:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 277:73]
  wire [22:0] _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 281:16]
  wire [22:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 280:12]
  wire [9:0] _io_out_T = {signOut,expOut}; // @[RoundAnyRawFNToRecFN.scala 286:23]
  assign io_out = {_io_out_T,fractOut}; // @[RoundAnyRawFNToRecFN.scala 286:33]
endmodule
module RoundRawFNToRecFN_e8_s24(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  output [32:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 310:15]
  RoundAnyRawFNToRecFN_ie8_is26_oe8_os24 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 310:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 318:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 315:44]
endmodule
module MulRecFN(
  input  [32:0] io_a,
  input  [32:0] io_b,
  output [32:0] io_out
);
  wire  mulRawFN__io_a_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_a_sExp; // @[MulRecFN.scala 113:26]
  wire [24:0] mulRawFN__io_a_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_b_sExp; // @[MulRecFN.scala 113:26]
  wire [24:0] mulRawFN__io_b_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_invalidExc; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 113:26]
  wire [9:0] mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 113:26]
  wire [26:0] mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 113:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulRecFN.scala 121:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[MulRecFN.scala 121:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[MulRecFN.scala 121:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[MulRecFN.scala 121:15]
  wire [8:0] mulRawFN_io_a_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  mulRawFN_io_a_isZero = mulRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  mulRawFN_io_a_isSpecial = mulRawFN_io_a_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _mulRawFN_io_a_out_sig_T = ~mulRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _mulRawFN_io_a_out_sig_T_1 = {1'h0,_mulRawFN_io_a_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  wire [8:0] mulRawFN_io_b_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  mulRawFN_io_b_isZero = mulRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  mulRawFN_io_b_isSpecial = mulRawFN_io_b_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _mulRawFN_io_b_out_sig_T = ~mulRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _mulRawFN_io_b_out_sig_T_1 = {1'h0,_mulRawFN_io_b_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  MulRawFN mulRawFN_ ( // @[MulRecFN.scala 113:26]
    .io_a_isNaN(mulRawFN__io_a_isNaN),
    .io_a_isInf(mulRawFN__io_a_isInf),
    .io_a_isZero(mulRawFN__io_a_isZero),
    .io_a_sign(mulRawFN__io_a_sign),
    .io_a_sExp(mulRawFN__io_a_sExp),
    .io_a_sig(mulRawFN__io_a_sig),
    .io_b_isNaN(mulRawFN__io_b_isNaN),
    .io_b_isInf(mulRawFN__io_b_isInf),
    .io_b_isZero(mulRawFN__io_b_isZero),
    .io_b_sign(mulRawFN__io_b_sign),
    .io_b_sExp(mulRawFN__io_b_sExp),
    .io_b_sig(mulRawFN__io_b_sig),
    .io_invalidExc(mulRawFN__io_invalidExc),
    .io_rawOut_isNaN(mulRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(mulRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(mulRawFN__io_rawOut_isZero),
    .io_rawOut_sign(mulRawFN__io_rawOut_sign),
    .io_rawOut_sExp(mulRawFN__io_rawOut_sExp),
    .io_rawOut_sig(mulRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN_e8_s24 roundRawFNToRecFN ( // @[MulRecFN.scala 121:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[MulRecFN.scala 127:23]
  assign mulRawFN__io_a_isNaN = mulRawFN_io_a_isSpecial & mulRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_a_isInf = mulRawFN_io_a_isSpecial & ~mulRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign mulRawFN__io_a_isZero = mulRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign mulRawFN__io_a_sign = io_a[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign mulRawFN__io_a_sExp = {1'b0,$signed(mulRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign mulRawFN__io_a_sig = {_mulRawFN_io_a_out_sig_T_1,io_a[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign mulRawFN__io_b_isNaN = mulRawFN_io_b_isSpecial & mulRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_b_isInf = mulRawFN_io_b_isSpecial & ~mulRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign mulRawFN__io_b_isZero = mulRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign mulRawFN__io_b_sign = io_b[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign mulRawFN__io_b_sExp = {1'b0,$signed(mulRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign mulRawFN__io_b_sig = {_mulRawFN_io_b_out_sig_T_1,io_b[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign roundRawFNToRecFN_io_invalidExc = mulRawFN__io_invalidExc; // @[MulRecFN.scala 122:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isInf = mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isZero = mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sign = mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sExp = mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sig = mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 124:39]
endmodule
module FP32Multiplier(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire [32:0] mulRecFN_io_a; // @[FPU.scala 88:26]
  wire [32:0] mulRecFN_io_b; // @[FPU.scala 88:26]
  wire [32:0] mulRecFN_io_out; // @[FPU.scala 88:26]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = mulRecFN_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = mulRecFN_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,mulRecFN_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  MulRecFN mulRecFN ( // @[FPU.scala 88:26]
    .io_a(mulRecFN_io_a),
    .io_b(mulRecFN_io_b),
    .io_out(mulRecFN_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign mulRecFN_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign mulRecFN_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module AddRawFN(
  input         io_subOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig
);
  wire  effSignB = io_b_sign ^ io_subOp; // @[AddRecFN.scala 60:30]
  wire  eqSigns = io_a_sign == effSignB; // @[AddRecFN.scala 61:29]
  wire [9:0] sDiffExps = $signed(io_a_sExp) - $signed(io_b_sExp); // @[AddRecFN.scala 63:31]
  wire  _modNatAlignDist_T = $signed(sDiffExps) < 10'sh0; // @[AddRecFN.scala 64:41]
  wire [9:0] _modNatAlignDist_T_3 = $signed(io_b_sExp) - $signed(io_a_sExp); // @[AddRecFN.scala 64:58]
  wire [9:0] _modNatAlignDist_T_4 = $signed(sDiffExps) < 10'sh0 ? $signed(_modNatAlignDist_T_3) : $signed(sDiffExps); // @[AddRecFN.scala 64:30]
  wire [4:0] modNatAlignDist = _modNatAlignDist_T_4[4:0]; // @[AddRecFN.scala 64:81]
  wire [4:0] _isMaxAlign_T = sDiffExps[9:5]; // @[AddRecFN.scala 66:19]
  wire  _isMaxAlign_T_6 = $signed(_isMaxAlign_T) != -5'sh1 | sDiffExps[4:0] == 5'h0; // @[AddRecFN.scala 67:51]
  wire  isMaxAlign = $signed(_isMaxAlign_T) != 5'sh0 & _isMaxAlign_T_6; // @[AddRecFN.scala 66:45]
  wire [4:0] alignDist = isMaxAlign ? 5'h1f : modNatAlignDist; // @[AddRecFN.scala 68:24]
  wire  _closeSubMags_T = ~eqSigns; // @[AddRecFN.scala 69:24]
  wire  closeSubMags = ~eqSigns & ~isMaxAlign & modNatAlignDist <= 5'h1; // @[AddRecFN.scala 69:48]
  wire  _close_alignedSigA_T = 10'sh0 <= $signed(sDiffExps); // @[AddRecFN.scala 73:18]
  wire [26:0] _close_alignedSigA_T_3 = {io_a_sig, 2'h0}; // @[AddRecFN.scala 73:58]
  wire [26:0] _close_alignedSigA_T_4 = 10'sh0 <= $signed(sDiffExps) & sDiffExps[0] ? _close_alignedSigA_T_3 : 27'h0; // @[AddRecFN.scala 73:12]
  wire [25:0] _close_alignedSigA_T_9 = {io_a_sig, 1'h0}; // @[AddRecFN.scala 74:58]
  wire [25:0] _close_alignedSigA_T_10 = _close_alignedSigA_T & ~sDiffExps[0] ? _close_alignedSigA_T_9 : 26'h0; // @[AddRecFN.scala 74:12]
  wire [26:0] _GEN_0 = {{1'd0}, _close_alignedSigA_T_10}; // @[AddRecFN.scala 73:68]
  wire [26:0] _close_alignedSigA_T_11 = _close_alignedSigA_T_4 | _GEN_0; // @[AddRecFN.scala 73:68]
  wire [24:0] _close_alignedSigA_T_13 = _modNatAlignDist_T ? io_a_sig : 25'h0; // @[AddRecFN.scala 75:12]
  wire [26:0] _GEN_1 = {{2'd0}, _close_alignedSigA_T_13}; // @[AddRecFN.scala 74:68]
  wire [26:0] _close_sSigSum_T = _close_alignedSigA_T_11 | _GEN_1; // @[AddRecFN.scala 76:43]
  wire [25:0] _close_sSigSum_T_2 = {io_b_sig, 1'h0}; // @[AddRecFN.scala 76:66]
  wire [26:0] _GEN_2 = {{1{_close_sSigSum_T_2[25]}},_close_sSigSum_T_2}; // @[AddRecFN.scala 76:50]
  wire [26:0] close_sSigSum = $signed(_close_sSigSum_T) - $signed(_GEN_2); // @[AddRecFN.scala 76:50]
  wire  _close_sigSum_T = $signed(close_sSigSum) < 27'sh0; // @[AddRecFN.scala 77:42]
  wire [26:0] _close_sigSum_T_3 = 27'sh0 - $signed(close_sSigSum); // @[AddRecFN.scala 77:49]
  wire [26:0] _close_sigSum_T_4 = $signed(close_sSigSum) < 27'sh0 ? $signed(_close_sigSum_T_3) : $signed(close_sSigSum); // @[AddRecFN.scala 77:27]
  wire [25:0] close_sigSum = _close_sigSum_T_4[25:0]; // @[AddRecFN.scala 77:79]
  wire  close_reduced2SigSum_reducedVec_0 = |close_sigSum[1:0]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_1 = |close_sigSum[3:2]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_2 = |close_sigSum[5:4]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_3 = |close_sigSum[7:6]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_4 = |close_sigSum[9:8]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_5 = |close_sigSum[11:10]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_6 = |close_sigSum[13:12]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_7 = |close_sigSum[15:14]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_8 = |close_sigSum[17:16]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_9 = |close_sigSum[19:18]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_10 = |close_sigSum[21:20]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_11 = |close_sigSum[23:22]; // @[primitives.scala 103:54]
  wire  close_reduced2SigSum_reducedVec_12 = |close_sigSum[25:24]; // @[primitives.scala 106:57]
  wire [5:0] close_reduced2SigSum_lo = {close_reduced2SigSum_reducedVec_5,close_reduced2SigSum_reducedVec_4,
    close_reduced2SigSum_reducedVec_3,close_reduced2SigSum_reducedVec_2,close_reduced2SigSum_reducedVec_1,
    close_reduced2SigSum_reducedVec_0}; // @[primitives.scala 107:20]
  wire [12:0] close_reduced2SigSum = {close_reduced2SigSum_reducedVec_12,close_reduced2SigSum_reducedVec_11,
    close_reduced2SigSum_reducedVec_10,close_reduced2SigSum_reducedVec_9,close_reduced2SigSum_reducedVec_8,
    close_reduced2SigSum_reducedVec_7,close_reduced2SigSum_reducedVec_6,close_reduced2SigSum_lo}; // @[primitives.scala 107:20]
  wire [3:0] _close_normDistReduced2_T_13 = close_reduced2SigSum[1] ? 4'hb : 4'hc; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_14 = close_reduced2SigSum[2] ? 4'ha : _close_normDistReduced2_T_13; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_15 = close_reduced2SigSum[3] ? 4'h9 : _close_normDistReduced2_T_14; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_16 = close_reduced2SigSum[4] ? 4'h8 : _close_normDistReduced2_T_15; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_17 = close_reduced2SigSum[5] ? 4'h7 : _close_normDistReduced2_T_16; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_18 = close_reduced2SigSum[6] ? 4'h6 : _close_normDistReduced2_T_17; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_19 = close_reduced2SigSum[7] ? 4'h5 : _close_normDistReduced2_T_18; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_20 = close_reduced2SigSum[8] ? 4'h4 : _close_normDistReduced2_T_19; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_21 = close_reduced2SigSum[9] ? 4'h3 : _close_normDistReduced2_T_20; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_22 = close_reduced2SigSum[10] ? 4'h2 : _close_normDistReduced2_T_21; // @[Mux.scala 47:70]
  wire [3:0] _close_normDistReduced2_T_23 = close_reduced2SigSum[11] ? 4'h1 : _close_normDistReduced2_T_22; // @[Mux.scala 47:70]
  wire [3:0] close_normDistReduced2 = close_reduced2SigSum[12] ? 4'h0 : _close_normDistReduced2_T_23; // @[Mux.scala 47:70]
  wire [4:0] close_nearNormDist = {close_normDistReduced2, 1'h0}; // @[AddRecFN.scala 81:53]
  wire [56:0] _GEN_7 = {{31'd0}, close_sigSum}; // @[AddRecFN.scala 82:38]
  wire [56:0] _close_sigOut_T = _GEN_7 << close_nearNormDist; // @[AddRecFN.scala 82:38]
  wire [57:0] _close_sigOut_T_1 = {_close_sigOut_T, 1'h0}; // @[AddRecFN.scala 82:59]
  wire [26:0] close_sigOut = _close_sigOut_T_1[26:0]; // @[AddRecFN.scala 82:63]
  wire  close_totalCancellation = ~(|close_sigOut[26:25]); // @[AddRecFN.scala 83:35]
  wire  close_notTotalCancellation_signOut = io_a_sign ^ _close_sigSum_T; // @[AddRecFN.scala 84:56]
  wire  far_signOut = _modNatAlignDist_T ? effSignB : io_a_sign; // @[AddRecFN.scala 87:26]
  wire [24:0] _far_sigLarger_T_1 = _modNatAlignDist_T ? io_b_sig : io_a_sig; // @[AddRecFN.scala 88:29]
  wire [23:0] far_sigLarger = _far_sigLarger_T_1[23:0]; // @[AddRecFN.scala 88:66]
  wire [24:0] _far_sigSmaller_T_1 = _modNatAlignDist_T ? io_a_sig : io_b_sig; // @[AddRecFN.scala 89:29]
  wire [23:0] far_sigSmaller = _far_sigSmaller_T_1[23:0]; // @[AddRecFN.scala 89:66]
  wire [28:0] _far_mainAlignedSigSmaller_T = {far_sigSmaller, 5'h0}; // @[AddRecFN.scala 90:52]
  wire [28:0] far_mainAlignedSigSmaller = _far_mainAlignedSigSmaller_T >> alignDist; // @[AddRecFN.scala 90:56]
  wire [25:0] _far_reduced4SigSmaller_T = {far_sigSmaller, 2'h0}; // @[AddRecFN.scala 91:60]
  wire  far_reduced4SigSmaller_reducedVec_0 = |_far_reduced4SigSmaller_T[3:0]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_1 = |_far_reduced4SigSmaller_T[7:4]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_2 = |_far_reduced4SigSmaller_T[11:8]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_3 = |_far_reduced4SigSmaller_T[15:12]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_4 = |_far_reduced4SigSmaller_T[19:16]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_5 = |_far_reduced4SigSmaller_T[23:20]; // @[primitives.scala 120:54]
  wire  far_reduced4SigSmaller_reducedVec_6 = |_far_reduced4SigSmaller_T[25:24]; // @[primitives.scala 123:57]
  wire [6:0] far_reduced4SigSmaller = {far_reduced4SigSmaller_reducedVec_6,far_reduced4SigSmaller_reducedVec_5,
    far_reduced4SigSmaller_reducedVec_4,far_reduced4SigSmaller_reducedVec_3,far_reduced4SigSmaller_reducedVec_2,
    far_reduced4SigSmaller_reducedVec_1,far_reduced4SigSmaller_reducedVec_0}; // @[primitives.scala 124:20]
  wire [8:0] far_roundExtraMask_shift = 9'sh100 >>> alignDist[4:2]; // @[primitives.scala 76:56]
  wire [6:0] far_roundExtraMask = {far_roundExtraMask_shift[1],far_roundExtraMask_shift[2],far_roundExtraMask_shift[3],
    far_roundExtraMask_shift[4],far_roundExtraMask_shift[5],far_roundExtraMask_shift[6],far_roundExtraMask_shift[7]}; // @[Cat.scala 33:92]
  wire [6:0] _far_alignedSigSmaller_T_3 = far_reduced4SigSmaller & far_roundExtraMask; // @[AddRecFN.scala 95:76]
  wire  _far_alignedSigSmaller_T_5 = |far_mainAlignedSigSmaller[2:0] | |_far_alignedSigSmaller_T_3; // @[AddRecFN.scala 95:49]
  wire [26:0] far_alignedSigSmaller = {far_mainAlignedSigSmaller[28:3],_far_alignedSigSmaller_T_5}; // @[Cat.scala 33:92]
  wire [26:0] _far_negAlignedSigSmaller_T = ~far_alignedSigSmaller; // @[AddRecFN.scala 97:62]
  wire [27:0] _far_negAlignedSigSmaller_T_1 = {1'h1,_far_negAlignedSigSmaller_T}; // @[Cat.scala 33:92]
  wire [27:0] far_negAlignedSigSmaller = _closeSubMags_T ? _far_negAlignedSigSmaller_T_1 : {{1'd0},
    far_alignedSigSmaller}; // @[AddRecFN.scala 97:39]
  wire [26:0] _far_sigSum_T = {far_sigLarger, 3'h0}; // @[AddRecFN.scala 98:36]
  wire [27:0] _GEN_3 = {{1'd0}, _far_sigSum_T}; // @[AddRecFN.scala 98:41]
  wire [27:0] _far_sigSum_T_2 = _GEN_3 + far_negAlignedSigSmaller; // @[AddRecFN.scala 98:41]
  wire [27:0] _GEN_4 = {{27'd0}, _closeSubMags_T}; // @[AddRecFN.scala 98:68]
  wire [27:0] far_sigSum = _far_sigSum_T_2 + _GEN_4; // @[AddRecFN.scala 98:68]
  wire [26:0] _GEN_5 = {{26'd0}, far_sigSum[0]}; // @[AddRecFN.scala 99:67]
  wire [26:0] _far_sigOut_T_2 = far_sigSum[27:1] | _GEN_5; // @[AddRecFN.scala 99:67]
  wire [27:0] _far_sigOut_T_3 = _closeSubMags_T ? far_sigSum : {{1'd0}, _far_sigOut_T_2}; // @[AddRecFN.scala 99:25]
  wire [26:0] far_sigOut = _far_sigOut_T_3[26:0]; // @[AddRecFN.scala 99:83]
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isInf & _closeSubMags_T; // @[AddRecFN.scala 102:57]
  wire  notNaN_isInfOut = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  wire  addZeros = io_a_isZero & io_b_isZero; // @[AddRecFN.scala 104:32]
  wire  notNaN_specialCase = notNaN_isInfOut | addZeros; // @[AddRecFN.scala 105:46]
  wire  _notNaN_signOut_T_1 = io_a_isInf & io_a_sign; // @[AddRecFN.scala 109:39]
  wire  _notNaN_signOut_T_2 = eqSigns & io_a_sign | _notNaN_signOut_T_1; // @[AddRecFN.scala 108:63]
  wire  _notNaN_signOut_T_3 = io_b_isInf & effSignB; // @[AddRecFN.scala 110:39]
  wire  _notNaN_signOut_T_4 = _notNaN_signOut_T_2 | _notNaN_signOut_T_3; // @[AddRecFN.scala 109:63]
  wire  _notNaN_signOut_T_9 = ~notNaN_specialCase; // @[AddRecFN.scala 112:10]
  wire  _notNaN_signOut_T_12 = ~notNaN_specialCase & closeSubMags & ~close_totalCancellation; // @[AddRecFN.scala 112:46]
  wire  _notNaN_signOut_T_13 = _notNaN_signOut_T_12 & close_notTotalCancellation_signOut; // @[AddRecFN.scala 113:38]
  wire  _notNaN_signOut_T_14 = _notNaN_signOut_T_4 | _notNaN_signOut_T_13; // @[AddRecFN.scala 111:63]
  wire  _notNaN_signOut_T_18 = _notNaN_signOut_T_9 & ~closeSubMags & far_signOut; // @[AddRecFN.scala 114:47]
  wire [9:0] _common_sExpOut_T_2 = closeSubMags | _modNatAlignDist_T ? $signed(io_b_sExp) : $signed(io_a_sExp); // @[AddRecFN.scala 116:13]
  wire [4:0] _common_sExpOut_T_3 = closeSubMags ? close_nearNormDist : {{4'd0}, _closeSubMags_T}; // @[AddRecFN.scala 117:18]
  wire [5:0] _common_sExpOut_T_4 = {1'b0,$signed(_common_sExpOut_T_3)}; // @[AddRecFN.scala 117:66]
  wire [9:0] _GEN_6 = {{4{_common_sExpOut_T_4[5]}},_common_sExpOut_T_4}; // @[AddRecFN.scala 117:13]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[AddRecFN.scala 121:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[AddRecFN.scala 125:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  assign io_rawOut_isZero = addZeros | ~notNaN_isInfOut & closeSubMags & close_totalCancellation; // @[AddRecFN.scala 106:37]
  assign io_rawOut_sign = _notNaN_signOut_T_14 | _notNaN_signOut_T_18; // @[AddRecFN.scala 113:77]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - $signed(_GEN_6); // @[AddRecFN.scala 117:13]
  assign io_rawOut_sig = closeSubMags ? close_sigOut : far_sigOut; // @[AddRecFN.scala 118:28]
endmodule
module AddRecFN(
  input         io_subOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  output [32:0] io_out
);
  wire  addRawFN__io_subOp; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_a_sExp; // @[AddRecFN.scala 147:26]
  wire [24:0] addRawFN__io_a_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_b_sExp; // @[AddRecFN.scala 147:26]
  wire [24:0] addRawFN__io_b_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_invalidExc; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_sign; // @[AddRecFN.scala 147:26]
  wire [9:0] addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 147:26]
  wire [26:0] addRawFN__io_rawOut_sig; // @[AddRecFN.scala 147:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[AddRecFN.scala 157:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[AddRecFN.scala 157:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[AddRecFN.scala 157:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[AddRecFN.scala 157:15]
  wire [8:0] addRawFN_io_a_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  addRawFN_io_a_isZero = addRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  addRawFN_io_a_isSpecial = addRawFN_io_a_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _addRawFN_io_a_out_sig_T = ~addRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _addRawFN_io_a_out_sig_T_1 = {1'h0,_addRawFN_io_a_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  wire [8:0] addRawFN_io_b_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  addRawFN_io_b_isZero = addRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  addRawFN_io_b_isSpecial = addRawFN_io_b_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _addRawFN_io_b_out_sig_T = ~addRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _addRawFN_io_b_out_sig_T_1 = {1'h0,_addRawFN_io_b_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  AddRawFN addRawFN_ ( // @[AddRecFN.scala 147:26]
    .io_subOp(addRawFN__io_subOp),
    .io_a_isNaN(addRawFN__io_a_isNaN),
    .io_a_isInf(addRawFN__io_a_isInf),
    .io_a_isZero(addRawFN__io_a_isZero),
    .io_a_sign(addRawFN__io_a_sign),
    .io_a_sExp(addRawFN__io_a_sExp),
    .io_a_sig(addRawFN__io_a_sig),
    .io_b_isNaN(addRawFN__io_b_isNaN),
    .io_b_isInf(addRawFN__io_b_isInf),
    .io_b_isZero(addRawFN__io_b_isZero),
    .io_b_sign(addRawFN__io_b_sign),
    .io_b_sExp(addRawFN__io_b_sExp),
    .io_b_sig(addRawFN__io_b_sig),
    .io_invalidExc(addRawFN__io_invalidExc),
    .io_rawOut_isNaN(addRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(addRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(addRawFN__io_rawOut_isZero),
    .io_rawOut_sign(addRawFN__io_rawOut_sign),
    .io_rawOut_sExp(addRawFN__io_rawOut_sExp),
    .io_rawOut_sig(addRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN_e8_s24 roundRawFNToRecFN ( // @[AddRecFN.scala 157:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[AddRecFN.scala 163:23]
  assign addRawFN__io_subOp = io_subOp; // @[AddRecFN.scala 149:30]
  assign addRawFN__io_a_isNaN = addRawFN_io_a_isSpecial & addRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_a_isInf = addRawFN_io_a_isSpecial & ~addRawFN_io_a_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign addRawFN__io_a_isZero = addRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign addRawFN__io_a_sign = io_a[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign addRawFN__io_a_sExp = {1'b0,$signed(addRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign addRawFN__io_a_sig = {_addRawFN_io_a_out_sig_T_1,io_a[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign addRawFN__io_b_isNaN = addRawFN_io_b_isSpecial & addRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_b_isInf = addRawFN_io_b_isSpecial & ~addRawFN_io_b_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  assign addRawFN__io_b_isZero = addRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign addRawFN__io_b_sign = io_b[32]; // @[rawFloatFromRecFN.scala 59:25]
  assign addRawFN__io_b_sExp = {1'b0,$signed(addRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign addRawFN__io_b_sig = {_addRawFN_io_b_out_sig_T_1,io_b[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign roundRawFNToRecFN_io_invalidExc = addRawFN__io_invalidExc; // @[AddRecFN.scala 158:39]
  assign roundRawFNToRecFN_io_in_isNaN = addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isInf = addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isZero = addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sign = addRawFN__io_rawOut_sign; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sExp = addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sig = addRawFN__io_rawOut_sig; // @[AddRecFN.scala 160:39]
endmodule
module FP32Sub(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire  adder_io_subOp; // @[FPU.scala 45:23]
  wire [32:0] adder_io_a; // @[FPU.scala 45:23]
  wire [32:0] adder_io_b; // @[FPU.scala 45:23]
  wire [32:0] adder_io_out; // @[FPU.scala 45:23]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = adder_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = adder_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,adder_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  AddRecFN adder ( // @[FPU.scala 45:23]
    .io_subOp(adder_io_subOp),
    .io_a(adder_io_a),
    .io_b(adder_io_b),
    .io_out(adder_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign adder_io_subOp = 1'h1; // @[FPU.scala 52:20]
  assign adder_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign adder_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module FP32Adder(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_result
);
  wire  adder_io_subOp; // @[FPU.scala 17:23]
  wire [32:0] adder_io_a; // @[FPU.scala 17:23]
  wire [32:0] adder_io_b; // @[FPU.scala 17:23]
  wire [32:0] adder_io_out; // @[FPU.scala 17:23]
  wire  a_recoded_rawIn_sign = io_a[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] a_recoded_rawIn_expIn = io_a[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] a_recoded_rawIn_fractIn = io_a[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  a_recoded_rawIn_isZeroExpIn = a_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  a_recoded_rawIn_isZeroFractIn = a_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _a_recoded_rawIn_normDist_T_23 = a_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_24 = a_recoded_rawIn_fractIn[2] ? 5'h14 : _a_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_25 = a_recoded_rawIn_fractIn[3] ? 5'h13 : _a_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_26 = a_recoded_rawIn_fractIn[4] ? 5'h12 : _a_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_27 = a_recoded_rawIn_fractIn[5] ? 5'h11 : _a_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_28 = a_recoded_rawIn_fractIn[6] ? 5'h10 : _a_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_29 = a_recoded_rawIn_fractIn[7] ? 5'hf : _a_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_30 = a_recoded_rawIn_fractIn[8] ? 5'he : _a_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_31 = a_recoded_rawIn_fractIn[9] ? 5'hd : _a_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_32 = a_recoded_rawIn_fractIn[10] ? 5'hc : _a_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_33 = a_recoded_rawIn_fractIn[11] ? 5'hb : _a_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_34 = a_recoded_rawIn_fractIn[12] ? 5'ha : _a_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_35 = a_recoded_rawIn_fractIn[13] ? 5'h9 : _a_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_36 = a_recoded_rawIn_fractIn[14] ? 5'h8 : _a_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_37 = a_recoded_rawIn_fractIn[15] ? 5'h7 : _a_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_38 = a_recoded_rawIn_fractIn[16] ? 5'h6 : _a_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_39 = a_recoded_rawIn_fractIn[17] ? 5'h5 : _a_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_40 = a_recoded_rawIn_fractIn[18] ? 5'h4 : _a_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_41 = a_recoded_rawIn_fractIn[19] ? 5'h3 : _a_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_42 = a_recoded_rawIn_fractIn[20] ? 5'h2 : _a_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _a_recoded_rawIn_normDist_T_43 = a_recoded_rawIn_fractIn[21] ? 5'h1 : _a_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] a_recoded_rawIn_normDist = a_recoded_rawIn_fractIn[22] ? 5'h0 : _a_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_8 = {{31'd0}, a_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _a_recoded_rawIn_subnormFract_T = _GEN_8 << a_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] a_recoded_rawIn_subnormFract = {_a_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_0 = {{4'd0}, a_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T = _GEN_0 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _a_recoded_rawIn_adjustedExp_T_1 = a_recoded_rawIn_isZeroExpIn ? _a_recoded_rawIn_adjustedExp_T : {{1'd0},
    a_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _a_recoded_rawIn_adjustedExp_T_2 = a_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_1 = {{6'd0}, _a_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _a_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_1; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_2 = {{1'd0}, _a_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] a_recoded_rawIn_adjustedExp = _a_recoded_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 57:9]
  wire  a_recoded_rawIn_isZero = a_recoded_rawIn_isZeroExpIn & a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  a_recoded_rawIn_isSpecial = a_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  a_recoded_rawIn__isNaN = a_recoded_rawIn_isSpecial & ~a_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] a_recoded_rawIn__sExp = {1'b0,$signed(a_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _a_recoded_rawIn_out_sig_T = ~a_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _a_recoded_rawIn_out_sig_T_2 = a_recoded_rawIn_isZeroExpIn ? a_recoded_rawIn_subnormFract :
    a_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] a_recoded_rawIn__sig = {1'h0,_a_recoded_rawIn_out_sig_T,_a_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _a_recoded_T_1 = a_recoded_rawIn_isZero ? 3'h0 : a_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_3 = {{2'd0}, a_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _a_recoded_T_3 = _a_recoded_T_1 | _GEN_3; // @[recFNFromFN.scala 48:76]
  wire [9:0] _a_recoded_T_6 = {a_recoded_rawIn_sign,_a_recoded_T_3,a_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire  b_recoded_rawIn_sign = io_b[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] b_recoded_rawIn_expIn = io_b[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] b_recoded_rawIn_fractIn = io_b[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  b_recoded_rawIn_isZeroExpIn = b_recoded_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  b_recoded_rawIn_isZeroFractIn = b_recoded_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _b_recoded_rawIn_normDist_T_23 = b_recoded_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_24 = b_recoded_rawIn_fractIn[2] ? 5'h14 : _b_recoded_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_25 = b_recoded_rawIn_fractIn[3] ? 5'h13 : _b_recoded_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_26 = b_recoded_rawIn_fractIn[4] ? 5'h12 : _b_recoded_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_27 = b_recoded_rawIn_fractIn[5] ? 5'h11 : _b_recoded_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_28 = b_recoded_rawIn_fractIn[6] ? 5'h10 : _b_recoded_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_29 = b_recoded_rawIn_fractIn[7] ? 5'hf : _b_recoded_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_30 = b_recoded_rawIn_fractIn[8] ? 5'he : _b_recoded_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_31 = b_recoded_rawIn_fractIn[9] ? 5'hd : _b_recoded_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_32 = b_recoded_rawIn_fractIn[10] ? 5'hc : _b_recoded_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_33 = b_recoded_rawIn_fractIn[11] ? 5'hb : _b_recoded_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_34 = b_recoded_rawIn_fractIn[12] ? 5'ha : _b_recoded_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_35 = b_recoded_rawIn_fractIn[13] ? 5'h9 : _b_recoded_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_36 = b_recoded_rawIn_fractIn[14] ? 5'h8 : _b_recoded_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_37 = b_recoded_rawIn_fractIn[15] ? 5'h7 : _b_recoded_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_38 = b_recoded_rawIn_fractIn[16] ? 5'h6 : _b_recoded_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_39 = b_recoded_rawIn_fractIn[17] ? 5'h5 : _b_recoded_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_40 = b_recoded_rawIn_fractIn[18] ? 5'h4 : _b_recoded_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_41 = b_recoded_rawIn_fractIn[19] ? 5'h3 : _b_recoded_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_42 = b_recoded_rawIn_fractIn[20] ? 5'h2 : _b_recoded_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _b_recoded_rawIn_normDist_T_43 = b_recoded_rawIn_fractIn[21] ? 5'h1 : _b_recoded_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] b_recoded_rawIn_normDist = b_recoded_rawIn_fractIn[22] ? 5'h0 : _b_recoded_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_9 = {{31'd0}, b_recoded_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _b_recoded_rawIn_subnormFract_T = _GEN_9 << b_recoded_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] b_recoded_rawIn_subnormFract = {_b_recoded_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_4 = {{4'd0}, b_recoded_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T = _GEN_4 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _b_recoded_rawIn_adjustedExp_T_1 = b_recoded_rawIn_isZeroExpIn ? _b_recoded_rawIn_adjustedExp_T : {{1'd0},
    b_recoded_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _b_recoded_rawIn_adjustedExp_T_2 = b_recoded_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_5 = {{6'd0}, _b_recoded_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _b_recoded_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_5; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_6 = {{1'd0}, _b_recoded_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] b_recoded_rawIn_adjustedExp = _b_recoded_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 57:9]
  wire  b_recoded_rawIn_isZero = b_recoded_rawIn_isZeroExpIn & b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  b_recoded_rawIn_isSpecial = b_recoded_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  b_recoded_rawIn__isNaN = b_recoded_rawIn_isSpecial & ~b_recoded_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] b_recoded_rawIn__sExp = {1'b0,$signed(b_recoded_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _b_recoded_rawIn_out_sig_T = ~b_recoded_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _b_recoded_rawIn_out_sig_T_2 = b_recoded_rawIn_isZeroExpIn ? b_recoded_rawIn_subnormFract :
    b_recoded_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] b_recoded_rawIn__sig = {1'h0,_b_recoded_rawIn_out_sig_T,_b_recoded_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _b_recoded_T_1 = b_recoded_rawIn_isZero ? 3'h0 : b_recoded_rawIn__sExp[8:6]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_7 = {{2'd0}, b_recoded_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _b_recoded_T_3 = _b_recoded_T_1 | _GEN_7; // @[recFNFromFN.scala 48:76]
  wire [9:0] _b_recoded_T_6 = {b_recoded_rawIn_sign,_b_recoded_T_3,b_recoded_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  wire [8:0] io_result_rawIn_exp = adder_io_out[31:23]; // @[rawFloatFromRecFN.scala 51:21]
  wire  io_result_rawIn_isZero = io_result_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  io_result_rawIn_isSpecial = io_result_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  io_result_rawIn__isNaN = io_result_rawIn_isSpecial & io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_result_rawIn__isInf = io_result_rawIn_isSpecial & ~io_result_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 57:33]
  wire  io_result_rawIn__sign = adder_io_out[32]; // @[rawFloatFromRecFN.scala 59:25]
  wire [9:0] io_result_rawIn__sExp = {1'b0,$signed(io_result_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _io_result_rawIn_out_sig_T = ~io_result_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [24:0] io_result_rawIn__sig = {1'h0,_io_result_rawIn_out_sig_T,adder_io_out[22:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  io_result_isSubnormal = $signed(io_result_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 51:38]
  wire [4:0] io_result_denormShiftDist = 5'h1 - io_result_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 52:35]
  wire [23:0] _io_result_denormFract_T_1 = io_result_rawIn__sig[24:1] >> io_result_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [22:0] io_result_denormFract = _io_result_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 53:60]
  wire [7:0] _io_result_expOut_T_2 = io_result_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 58:45]
  wire [7:0] _io_result_expOut_T_3 = io_result_isSubnormal ? 8'h0 : _io_result_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_result_expOut_T_4 = io_result_rawIn__isNaN | io_result_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [7:0] _io_result_expOut_T_6 = _io_result_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] io_result_expOut = _io_result_expOut_T_3 | _io_result_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [22:0] _io_result_fractOut_T_1 = io_result_rawIn__isInf ? 23'h0 : io_result_rawIn__sig[22:0]; // @[fNFromRecFN.scala 64:20]
  wire [22:0] io_result_fractOut = io_result_isSubnormal ? io_result_denormFract : _io_result_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [8:0] io_result_hi = {io_result_rawIn__sign,io_result_expOut}; // @[Cat.scala 33:92]
  AddRecFN adder ( // @[FPU.scala 17:23]
    .io_subOp(adder_io_subOp),
    .io_a(adder_io_a),
    .io_b(adder_io_b),
    .io_out(adder_io_out)
  );
  assign io_result = {io_result_hi,io_result_fractOut}; // @[Cat.scala 33:92]
  assign adder_io_subOp = 1'h0; // @[FPU.scala 24:20]
  assign adder_io_a = {_a_recoded_T_6,a_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  assign adder_io_b = {_b_recoded_T_6,b_recoded_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
endmodule
module FP32RoPEcore(
  input         clock,
  input         reset,
  input         io_EN,
  input  [31:0] io_x_0,
  input  [31:0] io_x_1,
  input  [31:0] io_sin,
  input  [31:0] io_cos,
  output [31:0] io_xhat_0,
  output [31:0] io_xhat_1,
  output        io_ENout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] FP32Mult0_io_a; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult0_io_b; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult0_io_result; // @[RoPEModuleFP32.scala 106:27]
  wire [31:0] FP32Mult1_io_a; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult1_io_b; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult1_io_result; // @[RoPEModuleFP32.scala 110:27]
  wire [31:0] FP32Mult2_io_a; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult2_io_b; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult2_io_result; // @[RoPEModuleFP32.scala 114:27]
  wire [31:0] FP32Mult3_io_a; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Mult3_io_b; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Mult3_io_result; // @[RoPEModuleFP32.scala 118:27]
  wire [31:0] FP32Sub_io_a; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32Sub_io_b; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32Sub_io_result; // @[RoPEModuleFP32.scala 131:25]
  wire [31:0] FP32add_io_a; // @[RoPEModuleFP32.scala 135:25]
  wire [31:0] FP32add_io_b; // @[RoPEModuleFP32.scala 135:25]
  wire [31:0] FP32add_io_result; // @[RoPEModuleFP32.scala 135:25]
  reg [31:0] stage1Reg_0; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_1; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_2; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage1Reg_3; // @[RoPEModuleFP32.scala 95:28]
  reg [31:0] stage2Reg_0; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_1; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_2; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage2Reg_3; // @[RoPEModuleFP32.scala 96:28]
  reg [31:0] stage3Reg_0; // @[RoPEModuleFP32.scala 97:28]
  reg [31:0] stage3Reg_1; // @[RoPEModuleFP32.scala 97:28]
  reg  enReg_0; // @[RoPEModuleFP32.scala 98:24]
  reg  enReg_1; // @[RoPEModuleFP32.scala 98:24]
  reg  enReg_2; // @[RoPEModuleFP32.scala 98:24]
  wire [31:0] _WIRE_1_0 = FP32Sub_io_result; // @[RoPEModuleFP32.scala 139:{25,25}]
  wire [31:0] _WIRE_1_1 = FP32add_io_result; // @[RoPEModuleFP32.scala 139:{25,25}]
  FP32Multiplier FP32Mult0 ( // @[RoPEModuleFP32.scala 106:27]
    .io_a(FP32Mult0_io_a),
    .io_b(FP32Mult0_io_b),
    .io_result(FP32Mult0_io_result)
  );
  FP32Multiplier FP32Mult1 ( // @[RoPEModuleFP32.scala 110:27]
    .io_a(FP32Mult1_io_a),
    .io_b(FP32Mult1_io_b),
    .io_result(FP32Mult1_io_result)
  );
  FP32Multiplier FP32Mult2 ( // @[RoPEModuleFP32.scala 114:27]
    .io_a(FP32Mult2_io_a),
    .io_b(FP32Mult2_io_b),
    .io_result(FP32Mult2_io_result)
  );
  FP32Multiplier FP32Mult3 ( // @[RoPEModuleFP32.scala 118:27]
    .io_a(FP32Mult3_io_a),
    .io_b(FP32Mult3_io_b),
    .io_result(FP32Mult3_io_result)
  );
  FP32Sub FP32Sub ( // @[RoPEModuleFP32.scala 131:25]
    .io_a(FP32Sub_io_a),
    .io_b(FP32Sub_io_b),
    .io_result(FP32Sub_io_result)
  );
  FP32Adder FP32add ( // @[RoPEModuleFP32.scala 135:25]
    .io_a(FP32add_io_a),
    .io_b(FP32add_io_b),
    .io_result(FP32add_io_result)
  );
  assign io_xhat_0 = enReg_2 ? stage3Reg_0 : 32'h0; // @[RoPEModuleFP32.scala 142:22]
  assign io_xhat_1 = enReg_2 ? stage3Reg_1 : 32'h0; // @[RoPEModuleFP32.scala 143:22]
  assign io_ENout = enReg_2; // @[RoPEModuleFP32.scala 144:14]
  assign FP32Mult0_io_a = stage1Reg_0; // @[RoPEModuleFP32.scala 107:20]
  assign FP32Mult0_io_b = stage1Reg_2; // @[RoPEModuleFP32.scala 108:20]
  assign FP32Mult1_io_a = stage1Reg_1; // @[RoPEModuleFP32.scala 111:20]
  assign FP32Mult1_io_b = stage1Reg_2; // @[RoPEModuleFP32.scala 112:20]
  assign FP32Mult2_io_a = stage1Reg_0; // @[RoPEModuleFP32.scala 115:20]
  assign FP32Mult2_io_b = stage1Reg_3; // @[RoPEModuleFP32.scala 116:20]
  assign FP32Mult3_io_a = stage1Reg_1; // @[RoPEModuleFP32.scala 119:20]
  assign FP32Mult3_io_b = stage1Reg_3; // @[RoPEModuleFP32.scala 120:20]
  assign FP32Sub_io_a = stage2Reg_2; // @[RoPEModuleFP32.scala 132:18]
  assign FP32Sub_io_b = stage2Reg_1; // @[RoPEModuleFP32.scala 133:18]
  assign FP32add_io_a = stage2Reg_3; // @[RoPEModuleFP32.scala 136:18]
  assign FP32add_io_b = stage2Reg_0; // @[RoPEModuleFP32.scala 137:18]
  always @(posedge clock) begin
    stage1Reg_0 <= io_x_0; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_1 <= io_x_1; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_2 <= io_sin; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage1Reg_3 <= io_cos; // @[RoPEModuleFP32.scala 95:{36,36}]
    stage2Reg_0 <= FP32Mult0_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_1 <= FP32Mult1_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_2 <= FP32Mult2_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    stage2Reg_3 <= FP32Mult3_io_result; // @[RoPEModuleFP32.scala 123:{25,25}]
    if (reset) begin // @[RoPEModuleFP32.scala 97:28]
      stage3Reg_0 <= 32'h0; // @[RoPEModuleFP32.scala 97:28]
    end else begin
      stage3Reg_0 <= _WIRE_1_0; // @[RoPEModuleFP32.scala 139:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 97:28]
      stage3Reg_1 <= 32'h0; // @[RoPEModuleFP32.scala 97:28]
    end else begin
      stage3Reg_1 <= _WIRE_1_1; // @[RoPEModuleFP32.scala 139:15]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_0 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_0 <= io_EN; // @[RoPEModuleFP32.scala 101:14]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_1 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_1 <= enReg_0; // @[RoPEModuleFP32.scala 102:14]
    end
    if (reset) begin // @[RoPEModuleFP32.scala 98:24]
      enReg_2 <= 1'h0; // @[RoPEModuleFP32.scala 98:24]
    end else begin
      enReg_2 <= enReg_1; // @[RoPEModuleFP32.scala 103:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage1Reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage1Reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stage1Reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stage2Reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stage2Reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stage2Reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage2Reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage3Reg_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage3Reg_1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  enReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  enReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  enReg_2 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multiLaneRoPEmoduleV2(
  input         clock,
  input         reset,
  input  [31:0] io_x_0_0,
  input  [31:0] io_x_0_1,
  input  [31:0] io_x_1_0,
  input  [31:0] io_x_1_1,
  input  [31:0] io_x_2_0,
  input  [31:0] io_x_2_1,
  input  [31:0] io_x_3_0,
  input  [31:0] io_x_3_1,
  input  [31:0] io_x_4_0,
  input  [31:0] io_x_4_1,
  input  [31:0] io_x_5_0,
  input  [31:0] io_x_5_1,
  input  [31:0] io_x_6_0,
  input  [31:0] io_x_6_1,
  input  [31:0] io_x_7_0,
  input  [31:0] io_x_7_1,
  input         io_EN,
  input  [31:0] io_m_0,
  input  [31:0] io_m_1,
  input  [31:0] io_m_2,
  input  [31:0] io_m_3,
  input  [31:0] io_m_4,
  input  [31:0] io_m_5,
  input  [31:0] io_m_6,
  input  [31:0] io_m_7,
  input  [31:0] io_baseIndex_0,
  input  [31:0] io_baseIndex_1,
  input  [31:0] io_baseIndex_2,
  input  [31:0] io_baseIndex_3,
  input  [31:0] io_baseIndex_4,
  input  [31:0] io_baseIndex_5,
  input  [31:0] io_baseIndex_6,
  input  [31:0] io_baseIndex_7,
  input  [31:0] io_ResMode_0,
  input  [31:0] io_ResMode_1,
  input  [31:0] io_ResMode_2,
  input  [31:0] io_ResMode_3,
  input  [31:0] io_ResMode_4,
  input  [31:0] io_ResMode_5,
  input  [31:0] io_ResMode_6,
  input  [31:0] io_ResMode_7,
  output [31:0] io_xhat_0_0,
  output [31:0] io_xhat_0_1,
  output [31:0] io_xhat_1_0,
  output [31:0] io_xhat_1_1,
  output [31:0] io_xhat_2_0,
  output [31:0] io_xhat_2_1,
  output [31:0] io_xhat_3_0,
  output [31:0] io_xhat_3_1,
  output [31:0] io_xhat_4_0,
  output [31:0] io_xhat_4_1,
  output [31:0] io_xhat_5_0,
  output [31:0] io_xhat_5_1,
  output [31:0] io_xhat_6_0,
  output [31:0] io_xhat_6_1,
  output [31:0] io_xhat_7_0,
  output [31:0] io_xhat_7_1,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
`endif // RANDOMIZE_REG_INIT
  wire  FP32radianCaclulatorV2_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_1_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_1_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_1_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_1_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_1_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_2_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_2_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_2_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_2_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_2_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_3_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_3_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_3_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_3_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_3_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_4_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_4_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_4_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_4_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_4_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_5_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_5_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_5_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_5_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_5_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_6_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_6_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_6_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_6_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_6_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_7_clock; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_7_reset; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_x_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_x_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_7_io_EN; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_m; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_baseIndex; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_ResMode; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_out; // @[RoPEModuleFP32v2.scala 47:15]
  wire  FP32radianCaclulatorV2_7_io_ENout; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_xFWD_0; // @[RoPEModuleFP32v2.scala 47:15]
  wire [31:0] FP32radianCaclulatorV2_7_io_xFWD_1; // @[RoPEModuleFP32v2.scala 47:15]
  wire  SinCosLut_clock; // @[RoPEModuleFP32v2.scala 49:27]
  wire  SinCosLut_reset; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_0_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_0_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_1_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_1_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_2_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_2_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_3_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_3_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_4_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_4_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_5_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_5_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_6_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_6_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_7_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_x_7_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire  SinCosLut_io_EN; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_2; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_3; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_4; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_5; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_6; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_angle_7; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_2; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_3; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_4; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_5; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_6; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_sinOut_7; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_2; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_3; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_4; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_5; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_6; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_cosOut_7; // @[RoPEModuleFP32v2.scala 49:27]
  wire  SinCosLut_io_ENout; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_0_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_0_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_1_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_1_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_2_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_2_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_3_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_3_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_4_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_4_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_5_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_5_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_6_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_6_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_7_0; // @[RoPEModuleFP32v2.scala 49:27]
  wire [31:0] SinCosLut_io_xFWD_7_1; // @[RoPEModuleFP32v2.scala 49:27]
  wire  FP32RoPEcore_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_1_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_1_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_1_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_1_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_1_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_2_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_2_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_2_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_2_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_2_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_3_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_3_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_3_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_3_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_3_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_4_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_4_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_4_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_4_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_4_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_5_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_5_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_5_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_5_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_5_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_6_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_6_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_6_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_6_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_6_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_7_clock; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_7_reset; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_7_io_EN; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_x_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_x_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_sin; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_cos; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_xhat_0; // @[RoPEModuleFP32v2.scala 51:15]
  wire [31:0] FP32RoPEcore_7_io_xhat_1; // @[RoPEModuleFP32v2.scala 51:15]
  wire  FP32RoPEcore_7_io_ENout; // @[RoPEModuleFP32v2.scala 51:15]
  reg [31:0] stage1Reg_0_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_0_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_0_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_0_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_0_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_1_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_1_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_1_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_1_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_1_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_2_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_2_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_2_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_2_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_2_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_3_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_3_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_3_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_3_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_3_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_4_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_4_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_4_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_4_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_4_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_5_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_5_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_5_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_5_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_5_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_6_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_6_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_6_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_6_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_6_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_7_0; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_7_1; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_7_2; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_7_3; // @[RoPEModuleFP32v2.scala 55:28]
  reg [31:0] stage1Reg_7_4; // @[RoPEModuleFP32v2.scala 55:28]
  reg  stage1EN; // @[RoPEModuleFP32v2.scala 56:28]
  reg [31:0] stage2Reg_0_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_0_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_0_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_1_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_1_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_1_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_2_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_2_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_2_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_3_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_3_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_3_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_4_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_4_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_4_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_5_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_5_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_5_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_6_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_6_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_6_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_7_0; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_7_1; // @[RoPEModuleFP32v2.scala 57:28]
  reg [31:0] stage2Reg_7_2; // @[RoPEModuleFP32v2.scala 57:28]
  reg  stage2EN; // @[RoPEModuleFP32v2.scala 58:28]
  reg [31:0] stage3Reg_0_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_0_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_0_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_0_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_1_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_1_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_1_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_1_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_2_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_2_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_2_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_2_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_3_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_3_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_3_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_3_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_4_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_4_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_4_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_4_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_5_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_5_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_5_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_5_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_6_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_6_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_6_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_6_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_7_0; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_7_1; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_7_2; // @[RoPEModuleFP32v2.scala 59:28]
  reg [31:0] stage3Reg_7_3; // @[RoPEModuleFP32v2.scala 59:28]
  reg  stage3EN; // @[RoPEModuleFP32v2.scala 60:28]
  reg [31:0] outputReg_0_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_0_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_1_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_1_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_2_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_2_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_3_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_3_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_4_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_4_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_5_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_5_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_6_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_6_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_7_0; // @[RoPEModuleFP32v2.scala 121:28]
  reg [31:0] outputReg_7_1; // @[RoPEModuleFP32v2.scala 121:28]
  reg  validReg; // @[RoPEModuleFP32v2.scala 122:27]
  FP32radianCaclulatorV2 FP32radianCaclulatorV2 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_clock),
    .reset(FP32radianCaclulatorV2_reset),
    .io_x_0(FP32radianCaclulatorV2_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_io_x_1),
    .io_EN(FP32radianCaclulatorV2_io_EN),
    .io_m(FP32radianCaclulatorV2_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_io_ResMode),
    .io_out(FP32radianCaclulatorV2_io_out),
    .io_ENout(FP32radianCaclulatorV2_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_1 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_1_clock),
    .reset(FP32radianCaclulatorV2_1_reset),
    .io_x_0(FP32radianCaclulatorV2_1_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_1_io_x_1),
    .io_EN(FP32radianCaclulatorV2_1_io_EN),
    .io_m(FP32radianCaclulatorV2_1_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_1_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_1_io_ResMode),
    .io_out(FP32radianCaclulatorV2_1_io_out),
    .io_ENout(FP32radianCaclulatorV2_1_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_1_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_1_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_2 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_2_clock),
    .reset(FP32radianCaclulatorV2_2_reset),
    .io_x_0(FP32radianCaclulatorV2_2_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_2_io_x_1),
    .io_EN(FP32radianCaclulatorV2_2_io_EN),
    .io_m(FP32radianCaclulatorV2_2_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_2_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_2_io_ResMode),
    .io_out(FP32radianCaclulatorV2_2_io_out),
    .io_ENout(FP32radianCaclulatorV2_2_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_2_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_2_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_3 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_3_clock),
    .reset(FP32radianCaclulatorV2_3_reset),
    .io_x_0(FP32radianCaclulatorV2_3_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_3_io_x_1),
    .io_EN(FP32radianCaclulatorV2_3_io_EN),
    .io_m(FP32radianCaclulatorV2_3_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_3_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_3_io_ResMode),
    .io_out(FP32radianCaclulatorV2_3_io_out),
    .io_ENout(FP32radianCaclulatorV2_3_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_3_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_3_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_4 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_4_clock),
    .reset(FP32radianCaclulatorV2_4_reset),
    .io_x_0(FP32radianCaclulatorV2_4_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_4_io_x_1),
    .io_EN(FP32radianCaclulatorV2_4_io_EN),
    .io_m(FP32radianCaclulatorV2_4_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_4_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_4_io_ResMode),
    .io_out(FP32radianCaclulatorV2_4_io_out),
    .io_ENout(FP32radianCaclulatorV2_4_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_4_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_4_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_5 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_5_clock),
    .reset(FP32radianCaclulatorV2_5_reset),
    .io_x_0(FP32radianCaclulatorV2_5_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_5_io_x_1),
    .io_EN(FP32radianCaclulatorV2_5_io_EN),
    .io_m(FP32radianCaclulatorV2_5_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_5_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_5_io_ResMode),
    .io_out(FP32radianCaclulatorV2_5_io_out),
    .io_ENout(FP32radianCaclulatorV2_5_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_5_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_5_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_6 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_6_clock),
    .reset(FP32radianCaclulatorV2_6_reset),
    .io_x_0(FP32radianCaclulatorV2_6_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_6_io_x_1),
    .io_EN(FP32radianCaclulatorV2_6_io_EN),
    .io_m(FP32radianCaclulatorV2_6_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_6_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_6_io_ResMode),
    .io_out(FP32radianCaclulatorV2_6_io_out),
    .io_ENout(FP32radianCaclulatorV2_6_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_6_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_6_io_xFWD_1)
  );
  FP32radianCaclulatorV2 FP32radianCaclulatorV2_7 ( // @[RoPEModuleFP32v2.scala 47:15]
    .clock(FP32radianCaclulatorV2_7_clock),
    .reset(FP32radianCaclulatorV2_7_reset),
    .io_x_0(FP32radianCaclulatorV2_7_io_x_0),
    .io_x_1(FP32radianCaclulatorV2_7_io_x_1),
    .io_EN(FP32radianCaclulatorV2_7_io_EN),
    .io_m(FP32radianCaclulatorV2_7_io_m),
    .io_baseIndex(FP32radianCaclulatorV2_7_io_baseIndex),
    .io_ResMode(FP32radianCaclulatorV2_7_io_ResMode),
    .io_out(FP32radianCaclulatorV2_7_io_out),
    .io_ENout(FP32radianCaclulatorV2_7_io_ENout),
    .io_xFWD_0(FP32radianCaclulatorV2_7_io_xFWD_0),
    .io_xFWD_1(FP32radianCaclulatorV2_7_io_xFWD_1)
  );
  multiPortSinCosModuleV2 SinCosLut ( // @[RoPEModuleFP32v2.scala 49:27]
    .clock(SinCosLut_clock),
    .reset(SinCosLut_reset),
    .io_x_0_0(SinCosLut_io_x_0_0),
    .io_x_0_1(SinCosLut_io_x_0_1),
    .io_x_1_0(SinCosLut_io_x_1_0),
    .io_x_1_1(SinCosLut_io_x_1_1),
    .io_x_2_0(SinCosLut_io_x_2_0),
    .io_x_2_1(SinCosLut_io_x_2_1),
    .io_x_3_0(SinCosLut_io_x_3_0),
    .io_x_3_1(SinCosLut_io_x_3_1),
    .io_x_4_0(SinCosLut_io_x_4_0),
    .io_x_4_1(SinCosLut_io_x_4_1),
    .io_x_5_0(SinCosLut_io_x_5_0),
    .io_x_5_1(SinCosLut_io_x_5_1),
    .io_x_6_0(SinCosLut_io_x_6_0),
    .io_x_6_1(SinCosLut_io_x_6_1),
    .io_x_7_0(SinCosLut_io_x_7_0),
    .io_x_7_1(SinCosLut_io_x_7_1),
    .io_EN(SinCosLut_io_EN),
    .io_angle_0(SinCosLut_io_angle_0),
    .io_angle_1(SinCosLut_io_angle_1),
    .io_angle_2(SinCosLut_io_angle_2),
    .io_angle_3(SinCosLut_io_angle_3),
    .io_angle_4(SinCosLut_io_angle_4),
    .io_angle_5(SinCosLut_io_angle_5),
    .io_angle_6(SinCosLut_io_angle_6),
    .io_angle_7(SinCosLut_io_angle_7),
    .io_sinOut_0(SinCosLut_io_sinOut_0),
    .io_sinOut_1(SinCosLut_io_sinOut_1),
    .io_sinOut_2(SinCosLut_io_sinOut_2),
    .io_sinOut_3(SinCosLut_io_sinOut_3),
    .io_sinOut_4(SinCosLut_io_sinOut_4),
    .io_sinOut_5(SinCosLut_io_sinOut_5),
    .io_sinOut_6(SinCosLut_io_sinOut_6),
    .io_sinOut_7(SinCosLut_io_sinOut_7),
    .io_cosOut_0(SinCosLut_io_cosOut_0),
    .io_cosOut_1(SinCosLut_io_cosOut_1),
    .io_cosOut_2(SinCosLut_io_cosOut_2),
    .io_cosOut_3(SinCosLut_io_cosOut_3),
    .io_cosOut_4(SinCosLut_io_cosOut_4),
    .io_cosOut_5(SinCosLut_io_cosOut_5),
    .io_cosOut_6(SinCosLut_io_cosOut_6),
    .io_cosOut_7(SinCosLut_io_cosOut_7),
    .io_ENout(SinCosLut_io_ENout),
    .io_xFWD_0_0(SinCosLut_io_xFWD_0_0),
    .io_xFWD_0_1(SinCosLut_io_xFWD_0_1),
    .io_xFWD_1_0(SinCosLut_io_xFWD_1_0),
    .io_xFWD_1_1(SinCosLut_io_xFWD_1_1),
    .io_xFWD_2_0(SinCosLut_io_xFWD_2_0),
    .io_xFWD_2_1(SinCosLut_io_xFWD_2_1),
    .io_xFWD_3_0(SinCosLut_io_xFWD_3_0),
    .io_xFWD_3_1(SinCosLut_io_xFWD_3_1),
    .io_xFWD_4_0(SinCosLut_io_xFWD_4_0),
    .io_xFWD_4_1(SinCosLut_io_xFWD_4_1),
    .io_xFWD_5_0(SinCosLut_io_xFWD_5_0),
    .io_xFWD_5_1(SinCosLut_io_xFWD_5_1),
    .io_xFWD_6_0(SinCosLut_io_xFWD_6_0),
    .io_xFWD_6_1(SinCosLut_io_xFWD_6_1),
    .io_xFWD_7_0(SinCosLut_io_xFWD_7_0),
    .io_xFWD_7_1(SinCosLut_io_xFWD_7_1)
  );
  FP32RoPEcore FP32RoPEcore ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_clock),
    .reset(FP32RoPEcore_reset),
    .io_EN(FP32RoPEcore_io_EN),
    .io_x_0(FP32RoPEcore_io_x_0),
    .io_x_1(FP32RoPEcore_io_x_1),
    .io_sin(FP32RoPEcore_io_sin),
    .io_cos(FP32RoPEcore_io_cos),
    .io_xhat_0(FP32RoPEcore_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_io_xhat_1),
    .io_ENout(FP32RoPEcore_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_1 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_1_clock),
    .reset(FP32RoPEcore_1_reset),
    .io_EN(FP32RoPEcore_1_io_EN),
    .io_x_0(FP32RoPEcore_1_io_x_0),
    .io_x_1(FP32RoPEcore_1_io_x_1),
    .io_sin(FP32RoPEcore_1_io_sin),
    .io_cos(FP32RoPEcore_1_io_cos),
    .io_xhat_0(FP32RoPEcore_1_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_1_io_xhat_1),
    .io_ENout(FP32RoPEcore_1_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_2 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_2_clock),
    .reset(FP32RoPEcore_2_reset),
    .io_EN(FP32RoPEcore_2_io_EN),
    .io_x_0(FP32RoPEcore_2_io_x_0),
    .io_x_1(FP32RoPEcore_2_io_x_1),
    .io_sin(FP32RoPEcore_2_io_sin),
    .io_cos(FP32RoPEcore_2_io_cos),
    .io_xhat_0(FP32RoPEcore_2_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_2_io_xhat_1),
    .io_ENout(FP32RoPEcore_2_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_3 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_3_clock),
    .reset(FP32RoPEcore_3_reset),
    .io_EN(FP32RoPEcore_3_io_EN),
    .io_x_0(FP32RoPEcore_3_io_x_0),
    .io_x_1(FP32RoPEcore_3_io_x_1),
    .io_sin(FP32RoPEcore_3_io_sin),
    .io_cos(FP32RoPEcore_3_io_cos),
    .io_xhat_0(FP32RoPEcore_3_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_3_io_xhat_1),
    .io_ENout(FP32RoPEcore_3_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_4 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_4_clock),
    .reset(FP32RoPEcore_4_reset),
    .io_EN(FP32RoPEcore_4_io_EN),
    .io_x_0(FP32RoPEcore_4_io_x_0),
    .io_x_1(FP32RoPEcore_4_io_x_1),
    .io_sin(FP32RoPEcore_4_io_sin),
    .io_cos(FP32RoPEcore_4_io_cos),
    .io_xhat_0(FP32RoPEcore_4_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_4_io_xhat_1),
    .io_ENout(FP32RoPEcore_4_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_5 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_5_clock),
    .reset(FP32RoPEcore_5_reset),
    .io_EN(FP32RoPEcore_5_io_EN),
    .io_x_0(FP32RoPEcore_5_io_x_0),
    .io_x_1(FP32RoPEcore_5_io_x_1),
    .io_sin(FP32RoPEcore_5_io_sin),
    .io_cos(FP32RoPEcore_5_io_cos),
    .io_xhat_0(FP32RoPEcore_5_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_5_io_xhat_1),
    .io_ENout(FP32RoPEcore_5_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_6 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_6_clock),
    .reset(FP32RoPEcore_6_reset),
    .io_EN(FP32RoPEcore_6_io_EN),
    .io_x_0(FP32RoPEcore_6_io_x_0),
    .io_x_1(FP32RoPEcore_6_io_x_1),
    .io_sin(FP32RoPEcore_6_io_sin),
    .io_cos(FP32RoPEcore_6_io_cos),
    .io_xhat_0(FP32RoPEcore_6_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_6_io_xhat_1),
    .io_ENout(FP32RoPEcore_6_io_ENout)
  );
  FP32RoPEcore FP32RoPEcore_7 ( // @[RoPEModuleFP32v2.scala 51:15]
    .clock(FP32RoPEcore_7_clock),
    .reset(FP32RoPEcore_7_reset),
    .io_EN(FP32RoPEcore_7_io_EN),
    .io_x_0(FP32RoPEcore_7_io_x_0),
    .io_x_1(FP32RoPEcore_7_io_x_1),
    .io_sin(FP32RoPEcore_7_io_sin),
    .io_cos(FP32RoPEcore_7_io_cos),
    .io_xhat_0(FP32RoPEcore_7_io_xhat_0),
    .io_xhat_1(FP32RoPEcore_7_io_xhat_1),
    .io_ENout(FP32RoPEcore_7_io_ENout)
  );
  assign io_xhat_0_0 = outputReg_0_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_0_1 = outputReg_0_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_1_0 = outputReg_1_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_1_1 = outputReg_1_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_2_0 = outputReg_2_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_2_1 = outputReg_2_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_3_0 = outputReg_3_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_3_1 = outputReg_3_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_4_0 = outputReg_4_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_4_1 = outputReg_4_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_5_0 = outputReg_5_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_5_1 = outputReg_5_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_6_0 = outputReg_6_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_6_1 = outputReg_6_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_xhat_7_0 = outputReg_7_0; // @[RoPEModuleFP32v2.scala 127:23]
  assign io_xhat_7_1 = outputReg_7_1; // @[RoPEModuleFP32v2.scala 128:23]
  assign io_valid = validReg; // @[RoPEModuleFP32v2.scala 130:14]
  assign FP32radianCaclulatorV2_clock = clock;
  assign FP32radianCaclulatorV2_reset = reset;
  assign FP32radianCaclulatorV2_io_x_0 = stage1Reg_0_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_io_x_1 = stage1Reg_0_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_io_m = stage1Reg_0_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_io_baseIndex = stage1Reg_0_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_io_ResMode = stage1Reg_0_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_1_clock = clock;
  assign FP32radianCaclulatorV2_1_reset = reset;
  assign FP32radianCaclulatorV2_1_io_x_0 = stage1Reg_1_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_1_io_x_1 = stage1Reg_1_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_1_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_1_io_m = stage1Reg_1_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_1_io_baseIndex = stage1Reg_1_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_1_io_ResMode = stage1Reg_1_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_2_clock = clock;
  assign FP32radianCaclulatorV2_2_reset = reset;
  assign FP32radianCaclulatorV2_2_io_x_0 = stage1Reg_2_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_2_io_x_1 = stage1Reg_2_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_2_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_2_io_m = stage1Reg_2_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_2_io_baseIndex = stage1Reg_2_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_2_io_ResMode = stage1Reg_2_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_3_clock = clock;
  assign FP32radianCaclulatorV2_3_reset = reset;
  assign FP32radianCaclulatorV2_3_io_x_0 = stage1Reg_3_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_3_io_x_1 = stage1Reg_3_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_3_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_3_io_m = stage1Reg_3_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_3_io_baseIndex = stage1Reg_3_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_3_io_ResMode = stage1Reg_3_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_4_clock = clock;
  assign FP32radianCaclulatorV2_4_reset = reset;
  assign FP32radianCaclulatorV2_4_io_x_0 = stage1Reg_4_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_4_io_x_1 = stage1Reg_4_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_4_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_4_io_m = stage1Reg_4_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_4_io_baseIndex = stage1Reg_4_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_4_io_ResMode = stage1Reg_4_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_5_clock = clock;
  assign FP32radianCaclulatorV2_5_reset = reset;
  assign FP32radianCaclulatorV2_5_io_x_0 = stage1Reg_5_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_5_io_x_1 = stage1Reg_5_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_5_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_5_io_m = stage1Reg_5_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_5_io_baseIndex = stage1Reg_5_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_5_io_ResMode = stage1Reg_5_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_6_clock = clock;
  assign FP32radianCaclulatorV2_6_reset = reset;
  assign FP32radianCaclulatorV2_6_io_x_0 = stage1Reg_6_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_6_io_x_1 = stage1Reg_6_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_6_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_6_io_m = stage1Reg_6_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_6_io_baseIndex = stage1Reg_6_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_6_io_ResMode = stage1Reg_6_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign FP32radianCaclulatorV2_7_clock = clock;
  assign FP32radianCaclulatorV2_7_reset = reset;
  assign FP32radianCaclulatorV2_7_io_x_0 = stage1Reg_7_0; // @[RoPEModuleFP32v2.scala 79:33]
  assign FP32radianCaclulatorV2_7_io_x_1 = stage1Reg_7_1; // @[RoPEModuleFP32v2.scala 80:33]
  assign FP32radianCaclulatorV2_7_io_EN = stage1EN; // @[RoPEModuleFP32v2.scala 78:33]
  assign FP32radianCaclulatorV2_7_io_m = stage1Reg_7_2; // @[RoPEModuleFP32v2.scala 81:33]
  assign FP32radianCaclulatorV2_7_io_baseIndex = stage1Reg_7_3; // @[RoPEModuleFP32v2.scala 82:33]
  assign FP32radianCaclulatorV2_7_io_ResMode = stage1Reg_7_4; // @[RoPEModuleFP32v2.scala 83:33]
  assign SinCosLut_clock = clock;
  assign SinCosLut_reset = reset;
  assign SinCosLut_io_x_0_0 = stage2Reg_0_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_0_1 = stage2Reg_0_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_1_0 = stage2Reg_1_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_1_1 = stage2Reg_1_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_2_0 = stage2Reg_2_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_2_1 = stage2Reg_2_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_3_0 = stage2Reg_3_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_3_1 = stage2Reg_3_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_4_0 = stage2Reg_4_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_4_1 = stage2Reg_4_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_5_0 = stage2Reg_5_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_5_1 = stage2Reg_5_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_6_0 = stage2Reg_6_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_6_1 = stage2Reg_6_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_x_7_0 = stage2Reg_7_0; // @[RoPEModuleFP32v2.scala 97:31]
  assign SinCosLut_io_x_7_1 = stage2Reg_7_1; // @[RoPEModuleFP32v2.scala 98:31]
  assign SinCosLut_io_EN = stage2EN; // @[RoPEModuleFP32v2.scala 95:21]
  assign SinCosLut_io_angle_0 = stage2Reg_0_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_1 = stage2Reg_1_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_2 = stage2Reg_2_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_3 = stage2Reg_3_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_4 = stage2Reg_4_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_5 = stage2Reg_5_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_6 = stage2Reg_6_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign SinCosLut_io_angle_7 = stage2Reg_7_2; // @[RoPEModuleFP32v2.scala 99:31]
  assign FP32RoPEcore_clock = clock;
  assign FP32RoPEcore_reset = reset;
  assign FP32RoPEcore_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_io_x_0 = stage3Reg_0_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_io_x_1 = stage3Reg_0_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_io_sin = stage3Reg_0_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_io_cos = stage3Reg_0_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_1_clock = clock;
  assign FP32RoPEcore_1_reset = reset;
  assign FP32RoPEcore_1_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_1_io_x_0 = stage3Reg_1_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_1_io_x_1 = stage3Reg_1_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_1_io_sin = stage3Reg_1_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_1_io_cos = stage3Reg_1_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_2_clock = clock;
  assign FP32RoPEcore_2_reset = reset;
  assign FP32RoPEcore_2_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_2_io_x_0 = stage3Reg_2_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_2_io_x_1 = stage3Reg_2_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_2_io_sin = stage3Reg_2_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_2_io_cos = stage3Reg_2_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_3_clock = clock;
  assign FP32RoPEcore_3_reset = reset;
  assign FP32RoPEcore_3_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_3_io_x_0 = stage3Reg_3_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_3_io_x_1 = stage3Reg_3_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_3_io_sin = stage3Reg_3_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_3_io_cos = stage3Reg_3_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_4_clock = clock;
  assign FP32RoPEcore_4_reset = reset;
  assign FP32RoPEcore_4_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_4_io_x_0 = stage3Reg_4_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_4_io_x_1 = stage3Reg_4_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_4_io_sin = stage3Reg_4_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_4_io_cos = stage3Reg_4_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_5_clock = clock;
  assign FP32RoPEcore_5_reset = reset;
  assign FP32RoPEcore_5_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_5_io_x_0 = stage3Reg_5_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_5_io_x_1 = stage3Reg_5_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_5_io_sin = stage3Reg_5_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_5_io_cos = stage3Reg_5_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_6_clock = clock;
  assign FP32RoPEcore_6_reset = reset;
  assign FP32RoPEcore_6_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_6_io_x_0 = stage3Reg_6_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_6_io_x_1 = stage3Reg_6_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_6_io_sin = stage3Reg_6_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_6_io_cos = stage3Reg_6_3; // @[RoPEModuleFP32v2.scala 117:29]
  assign FP32RoPEcore_7_clock = clock;
  assign FP32RoPEcore_7_reset = reset;
  assign FP32RoPEcore_7_io_EN = stage3EN; // @[RoPEModuleFP32v2.scala 113:29]
  assign FP32RoPEcore_7_io_x_0 = stage3Reg_7_0; // @[RoPEModuleFP32v2.scala 114:29]
  assign FP32RoPEcore_7_io_x_1 = stage3Reg_7_1; // @[RoPEModuleFP32v2.scala 115:29]
  assign FP32RoPEcore_7_io_sin = stage3Reg_7_2; // @[RoPEModuleFP32v2.scala 116:29]
  assign FP32RoPEcore_7_io_cos = stage3Reg_7_3; // @[RoPEModuleFP32v2.scala 117:29]
  always @(posedge clock) begin
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_0_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_0_0 <= io_x_0_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_0_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_0_1 <= io_x_0_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_0_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_0_2 <= io_m_0; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_0_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_0_3 <= io_baseIndex_0; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_0_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_0_4 <= io_ResMode_0; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_1_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_1_0 <= io_x_1_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_1_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_1_1 <= io_x_1_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_1_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_1_2 <= io_m_1; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_1_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_1_3 <= io_baseIndex_1; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_1_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_1_4 <= io_ResMode_1; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_2_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_2_0 <= io_x_2_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_2_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_2_1 <= io_x_2_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_2_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_2_2 <= io_m_2; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_2_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_2_3 <= io_baseIndex_2; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_2_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_2_4 <= io_ResMode_2; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_3_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_3_0 <= io_x_3_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_3_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_3_1 <= io_x_3_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_3_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_3_2 <= io_m_3; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_3_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_3_3 <= io_baseIndex_3; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_3_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_3_4 <= io_ResMode_3; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_4_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_4_0 <= io_x_4_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_4_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_4_1 <= io_x_4_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_4_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_4_2 <= io_m_4; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_4_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_4_3 <= io_baseIndex_4; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_4_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_4_4 <= io_ResMode_4; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_5_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_5_0 <= io_x_5_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_5_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_5_1 <= io_x_5_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_5_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_5_2 <= io_m_5; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_5_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_5_3 <= io_baseIndex_5; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_5_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_5_4 <= io_ResMode_5; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_6_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_6_0 <= io_x_6_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_6_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_6_1 <= io_x_6_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_6_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_6_2 <= io_m_6; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_6_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_6_3 <= io_baseIndex_6; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_6_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_6_4 <= io_ResMode_6; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_7_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_7_0 <= io_x_7_0; // @[RoPEModuleFP32v2.scala 65:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_7_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_7_1 <= io_x_7_1; // @[RoPEModuleFP32v2.scala 66:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_7_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_7_2 <= io_m_7; // @[RoPEModuleFP32v2.scala 67:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_7_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_7_3 <= io_baseIndex_7; // @[RoPEModuleFP32v2.scala 68:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 55:28]
      stage1Reg_7_4 <= 32'h0; // @[RoPEModuleFP32v2.scala 55:28]
    end else if (io_EN) begin // @[RoPEModuleFP32v2.scala 63:17]
      stage1Reg_7_4 <= io_ResMode_7; // @[RoPEModuleFP32v2.scala 69:29]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 56:28]
      stage1EN <= 1'h0; // @[RoPEModuleFP32v2.scala 56:28]
    end else begin
      stage1EN <= io_EN;
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_0_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_0_0 <= FP32radianCaclulatorV2_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_0_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_0_1 <= FP32radianCaclulatorV2_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_0_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_0_2 <= FP32radianCaclulatorV2_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_1_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_1_0 <= FP32radianCaclulatorV2_1_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_1_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_1_1 <= FP32radianCaclulatorV2_1_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_1_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_1_2 <= FP32radianCaclulatorV2_1_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_2_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_2_0 <= FP32radianCaclulatorV2_2_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_2_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_2_1 <= FP32radianCaclulatorV2_2_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_2_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_2_2 <= FP32radianCaclulatorV2_2_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_3_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_3_0 <= FP32radianCaclulatorV2_3_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_3_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_3_1 <= FP32radianCaclulatorV2_3_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_3_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_3_2 <= FP32radianCaclulatorV2_3_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_4_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_4_0 <= FP32radianCaclulatorV2_4_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_4_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_4_1 <= FP32radianCaclulatorV2_4_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_4_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_4_2 <= FP32radianCaclulatorV2_4_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_5_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_5_0 <= FP32radianCaclulatorV2_5_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_5_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_5_1 <= FP32radianCaclulatorV2_5_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_5_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_5_2 <= FP32radianCaclulatorV2_5_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_6_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_6_0 <= FP32radianCaclulatorV2_6_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_6_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_6_1 <= FP32radianCaclulatorV2_6_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_6_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_6_2 <= FP32radianCaclulatorV2_6_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_7_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_7_0 <= FP32radianCaclulatorV2_7_io_xFWD_0; // @[RoPEModuleFP32v2.scala 88:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_7_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_7_1 <= FP32radianCaclulatorV2_7_io_xFWD_1; // @[RoPEModuleFP32v2.scala 89:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 57:28]
      stage2Reg_7_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 57:28]
    end else begin
      stage2Reg_7_2 <= FP32radianCaclulatorV2_7_io_out; // @[RoPEModuleFP32v2.scala 90:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 58:28]
      stage2EN <= 1'h0; // @[RoPEModuleFP32v2.scala 58:28]
    end else begin
      stage2EN <= FP32radianCaclulatorV2_io_ENout; // @[RoPEModuleFP32v2.scala 92:14]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_0_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_0_0 <= SinCosLut_io_xFWD_0_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_0_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_0_1 <= SinCosLut_io_xFWD_0_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_0_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_0_2 <= SinCosLut_io_sinOut_0; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_0_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_0_3 <= SinCosLut_io_cosOut_0; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_1_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_1_0 <= SinCosLut_io_xFWD_1_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_1_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_1_1 <= SinCosLut_io_xFWD_1_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_1_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_1_2 <= SinCosLut_io_sinOut_1; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_1_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_1_3 <= SinCosLut_io_cosOut_1; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_2_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_2_0 <= SinCosLut_io_xFWD_2_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_2_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_2_1 <= SinCosLut_io_xFWD_2_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_2_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_2_2 <= SinCosLut_io_sinOut_2; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_2_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_2_3 <= SinCosLut_io_cosOut_2; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_3_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_3_0 <= SinCosLut_io_xFWD_3_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_3_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_3_1 <= SinCosLut_io_xFWD_3_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_3_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_3_2 <= SinCosLut_io_sinOut_3; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_3_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_3_3 <= SinCosLut_io_cosOut_3; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_4_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_4_0 <= SinCosLut_io_xFWD_4_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_4_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_4_1 <= SinCosLut_io_xFWD_4_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_4_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_4_2 <= SinCosLut_io_sinOut_4; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_4_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_4_3 <= SinCosLut_io_cosOut_4; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_5_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_5_0 <= SinCosLut_io_xFWD_5_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_5_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_5_1 <= SinCosLut_io_xFWD_5_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_5_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_5_2 <= SinCosLut_io_sinOut_5; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_5_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_5_3 <= SinCosLut_io_cosOut_5; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_6_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_6_0 <= SinCosLut_io_xFWD_6_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_6_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_6_1 <= SinCosLut_io_xFWD_6_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_6_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_6_2 <= SinCosLut_io_sinOut_6; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_6_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_6_3 <= SinCosLut_io_cosOut_6; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_7_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_7_0 <= SinCosLut_io_xFWD_7_0; // @[RoPEModuleFP32v2.scala 104:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_7_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_7_1 <= SinCosLut_io_xFWD_7_1; // @[RoPEModuleFP32v2.scala 105:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_7_2 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_7_2 <= SinCosLut_io_sinOut_7; // @[RoPEModuleFP32v2.scala 106:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 59:28]
      stage3Reg_7_3 <= 32'h0; // @[RoPEModuleFP32v2.scala 59:28]
    end else begin
      stage3Reg_7_3 <= SinCosLut_io_cosOut_7; // @[RoPEModuleFP32v2.scala 107:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 60:28]
      stage3EN <= 1'h0; // @[RoPEModuleFP32v2.scala 60:28]
    end else begin
      stage3EN <= SinCosLut_io_ENout; // @[RoPEModuleFP32v2.scala 109:14]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_0_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_0_0 <= FP32RoPEcore_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_0_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_0_1 <= FP32RoPEcore_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_1_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_1_0 <= FP32RoPEcore_1_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_1_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_1_1 <= FP32RoPEcore_1_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_2_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_2_0 <= FP32RoPEcore_2_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_2_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_2_1 <= FP32RoPEcore_2_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_3_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_3_0 <= FP32RoPEcore_3_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_3_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_3_1 <= FP32RoPEcore_3_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_4_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_4_0 <= FP32RoPEcore_4_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_4_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_4_1 <= FP32RoPEcore_4_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_5_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_5_0 <= FP32RoPEcore_5_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_5_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_5_1 <= FP32RoPEcore_5_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_6_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_6_0 <= FP32RoPEcore_6_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_6_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_6_1 <= FP32RoPEcore_6_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_7_0 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_7_0 <= FP32RoPEcore_7_io_xhat_0; // @[RoPEModuleFP32v2.scala 125:25]
    end
    if (reset) begin // @[RoPEModuleFP32v2.scala 121:28]
      outputReg_7_1 <= 32'h0; // @[RoPEModuleFP32v2.scala 121:28]
    end else begin
      outputReg_7_1 <= FP32RoPEcore_7_io_xhat_1; // @[RoPEModuleFP32v2.scala 126:25]
    end
    validReg <= FP32RoPEcore_io_ENout; // @[RoPEModuleFP32v2.scala 122:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage1Reg_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stage1Reg_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  stage1Reg_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  stage1Reg_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  stage1Reg_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  stage1Reg_1_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stage1Reg_1_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage1Reg_1_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage1Reg_1_3 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage1Reg_1_4 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stage1Reg_2_0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stage1Reg_2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stage1Reg_2_2 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  stage1Reg_2_3 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stage1Reg_2_4 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stage1Reg_3_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  stage1Reg_3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  stage1Reg_3_2 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  stage1Reg_3_3 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  stage1Reg_3_4 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stage1Reg_4_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stage1Reg_4_1 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stage1Reg_4_2 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  stage1Reg_4_3 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  stage1Reg_4_4 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  stage1Reg_5_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  stage1Reg_5_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  stage1Reg_5_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  stage1Reg_5_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  stage1Reg_5_4 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  stage1Reg_6_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  stage1Reg_6_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  stage1Reg_6_2 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  stage1Reg_6_3 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  stage1Reg_6_4 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  stage1Reg_7_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  stage1Reg_7_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  stage1Reg_7_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  stage1Reg_7_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  stage1Reg_7_4 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  stage1EN = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  stage2Reg_0_0 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  stage2Reg_0_1 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  stage2Reg_0_2 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  stage2Reg_1_0 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  stage2Reg_1_1 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  stage2Reg_1_2 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  stage2Reg_2_0 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  stage2Reg_2_1 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  stage2Reg_2_2 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  stage2Reg_3_0 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  stage2Reg_3_1 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  stage2Reg_3_2 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  stage2Reg_4_0 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  stage2Reg_4_1 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  stage2Reg_4_2 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  stage2Reg_5_0 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  stage2Reg_5_1 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  stage2Reg_5_2 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  stage2Reg_6_0 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  stage2Reg_6_1 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  stage2Reg_6_2 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  stage2Reg_7_0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  stage2Reg_7_1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  stage2Reg_7_2 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  stage2EN = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  stage3Reg_0_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  stage3Reg_0_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  stage3Reg_0_2 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  stage3Reg_0_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  stage3Reg_1_0 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  stage3Reg_1_1 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  stage3Reg_1_2 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  stage3Reg_1_3 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  stage3Reg_2_0 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  stage3Reg_2_1 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  stage3Reg_2_2 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  stage3Reg_2_3 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  stage3Reg_3_0 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  stage3Reg_3_1 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  stage3Reg_3_2 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  stage3Reg_3_3 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  stage3Reg_4_0 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  stage3Reg_4_1 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  stage3Reg_4_2 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  stage3Reg_4_3 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  stage3Reg_5_0 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  stage3Reg_5_1 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  stage3Reg_5_2 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  stage3Reg_5_3 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  stage3Reg_6_0 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  stage3Reg_6_1 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  stage3Reg_6_2 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  stage3Reg_6_3 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  stage3Reg_7_0 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  stage3Reg_7_1 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  stage3Reg_7_2 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  stage3Reg_7_3 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  stage3EN = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  outputReg_0_0 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  outputReg_0_1 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  outputReg_1_0 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  outputReg_1_1 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  outputReg_2_0 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  outputReg_2_1 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  outputReg_3_0 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  outputReg_3_1 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  outputReg_4_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  outputReg_4_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  outputReg_5_0 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  outputReg_5_1 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  outputReg_6_0 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  outputReg_6_1 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  outputReg_7_0 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  outputReg_7_1 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  validReg = _RAND_115[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
